VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiply_add_64x64
  CLASS BLOCK ;
  FOREIGN multiply_add_64x64 ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 27.570 10.640 30.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 10.640 210.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 10.640 390.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 10.640 570.670 688.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 688.400 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 92.520 700.000 93.120 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 133.320 700.000 133.920 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 137.400 700.000 138.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 141.480 700.000 142.080 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 145.560 700.000 146.160 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 149.640 700.000 150.240 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 153.720 700.000 154.320 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 157.800 700.000 158.400 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 161.880 700.000 162.480 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 165.960 700.000 166.560 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 170.040 700.000 170.640 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 96.600 700.000 97.200 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 174.120 700.000 174.720 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 178.200 700.000 178.800 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 182.280 700.000 182.880 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 186.360 700.000 186.960 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 190.440 700.000 191.040 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 194.520 700.000 195.120 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 198.600 700.000 199.200 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 202.680 700.000 203.280 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 206.760 700.000 207.360 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 210.840 700.000 211.440 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 100.680 700.000 101.280 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 214.920 700.000 215.520 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 219.000 700.000 219.600 ;
    END
  END a[31]
  PIN a[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 223.080 700.000 223.680 ;
    END
  END a[32]
  PIN a[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 227.160 700.000 227.760 ;
    END
  END a[33]
  PIN a[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.240 700.000 231.840 ;
    END
  END a[34]
  PIN a[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 235.320 700.000 235.920 ;
    END
  END a[35]
  PIN a[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 239.400 700.000 240.000 ;
    END
  END a[36]
  PIN a[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 243.480 700.000 244.080 ;
    END
  END a[37]
  PIN a[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 247.560 700.000 248.160 ;
    END
  END a[38]
  PIN a[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 251.640 700.000 252.240 ;
    END
  END a[39]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 104.760 700.000 105.360 ;
    END
  END a[3]
  PIN a[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 255.720 700.000 256.320 ;
    END
  END a[40]
  PIN a[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 259.800 700.000 260.400 ;
    END
  END a[41]
  PIN a[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 263.880 700.000 264.480 ;
    END
  END a[42]
  PIN a[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 267.960 700.000 268.560 ;
    END
  END a[43]
  PIN a[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 272.040 700.000 272.640 ;
    END
  END a[44]
  PIN a[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 276.120 700.000 276.720 ;
    END
  END a[45]
  PIN a[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 280.200 700.000 280.800 ;
    END
  END a[46]
  PIN a[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 284.280 700.000 284.880 ;
    END
  END a[47]
  PIN a[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 288.360 700.000 288.960 ;
    END
  END a[48]
  PIN a[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 292.440 700.000 293.040 ;
    END
  END a[49]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 108.840 700.000 109.440 ;
    END
  END a[4]
  PIN a[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 296.520 700.000 297.120 ;
    END
  END a[50]
  PIN a[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 300.600 700.000 301.200 ;
    END
  END a[51]
  PIN a[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 304.680 700.000 305.280 ;
    END
  END a[52]
  PIN a[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 308.760 700.000 309.360 ;
    END
  END a[53]
  PIN a[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 312.840 700.000 313.440 ;
    END
  END a[54]
  PIN a[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 316.920 700.000 317.520 ;
    END
  END a[55]
  PIN a[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 321.000 700.000 321.600 ;
    END
  END a[56]
  PIN a[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 325.080 700.000 325.680 ;
    END
  END a[57]
  PIN a[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 329.160 700.000 329.760 ;
    END
  END a[58]
  PIN a[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 333.240 700.000 333.840 ;
    END
  END a[59]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 112.920 700.000 113.520 ;
    END
  END a[5]
  PIN a[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 337.320 700.000 337.920 ;
    END
  END a[60]
  PIN a[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 341.400 700.000 342.000 ;
    END
  END a[61]
  PIN a[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 345.480 700.000 346.080 ;
    END
  END a[62]
  PIN a[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 349.560 700.000 350.160 ;
    END
  END a[63]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 117.000 700.000 117.600 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 121.080 700.000 121.680 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 125.160 700.000 125.760 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 129.240 700.000 129.840 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 353.640 700.000 354.240 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 394.440 700.000 395.040 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 398.520 700.000 399.120 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 402.600 700.000 403.200 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 406.680 700.000 407.280 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 410.760 700.000 411.360 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 414.840 700.000 415.440 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 418.920 700.000 419.520 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 423.000 700.000 423.600 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 427.080 700.000 427.680 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 431.160 700.000 431.760 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 357.720 700.000 358.320 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 435.240 700.000 435.840 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 439.320 700.000 439.920 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 443.400 700.000 444.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 447.480 700.000 448.080 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 451.560 700.000 452.160 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 455.640 700.000 456.240 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 459.720 700.000 460.320 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 463.800 700.000 464.400 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 467.880 700.000 468.480 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 471.960 700.000 472.560 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 361.800 700.000 362.400 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 476.040 700.000 476.640 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 480.120 700.000 480.720 ;
    END
  END b[31]
  PIN b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 484.200 700.000 484.800 ;
    END
  END b[32]
  PIN b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 488.280 700.000 488.880 ;
    END
  END b[33]
  PIN b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 492.360 700.000 492.960 ;
    END
  END b[34]
  PIN b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 496.440 700.000 497.040 ;
    END
  END b[35]
  PIN b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 500.520 700.000 501.120 ;
    END
  END b[36]
  PIN b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 504.600 700.000 505.200 ;
    END
  END b[37]
  PIN b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 508.680 700.000 509.280 ;
    END
  END b[38]
  PIN b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 512.760 700.000 513.360 ;
    END
  END b[39]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 365.880 700.000 366.480 ;
    END
  END b[3]
  PIN b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 516.840 700.000 517.440 ;
    END
  END b[40]
  PIN b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 520.920 700.000 521.520 ;
    END
  END b[41]
  PIN b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 525.000 700.000 525.600 ;
    END
  END b[42]
  PIN b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 529.080 700.000 529.680 ;
    END
  END b[43]
  PIN b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 533.160 700.000 533.760 ;
    END
  END b[44]
  PIN b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 537.240 700.000 537.840 ;
    END
  END b[45]
  PIN b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 541.320 700.000 541.920 ;
    END
  END b[46]
  PIN b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 545.400 700.000 546.000 ;
    END
  END b[47]
  PIN b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 549.480 700.000 550.080 ;
    END
  END b[48]
  PIN b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 553.560 700.000 554.160 ;
    END
  END b[49]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 369.960 700.000 370.560 ;
    END
  END b[4]
  PIN b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 557.640 700.000 558.240 ;
    END
  END b[50]
  PIN b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 561.720 700.000 562.320 ;
    END
  END b[51]
  PIN b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 565.800 700.000 566.400 ;
    END
  END b[52]
  PIN b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 569.880 700.000 570.480 ;
    END
  END b[53]
  PIN b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 573.960 700.000 574.560 ;
    END
  END b[54]
  PIN b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 578.040 700.000 578.640 ;
    END
  END b[55]
  PIN b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 582.120 700.000 582.720 ;
    END
  END b[56]
  PIN b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 586.200 700.000 586.800 ;
    END
  END b[57]
  PIN b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 590.280 700.000 590.880 ;
    END
  END b[58]
  PIN b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 594.360 700.000 594.960 ;
    END
  END b[59]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 374.040 700.000 374.640 ;
    END
  END b[5]
  PIN b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 598.440 700.000 599.040 ;
    END
  END b[60]
  PIN b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 602.520 700.000 603.120 ;
    END
  END b[61]
  PIN b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 606.600 700.000 607.200 ;
    END
  END b[62]
  PIN b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 610.680 700.000 611.280 ;
    END
  END b[63]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 378.120 700.000 378.720 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 382.200 700.000 382.800 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 386.280 700.000 386.880 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 696.000 390.360 700.000 390.960 ;
    END
  END b[9]
  PIN c[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END c[0]
  PIN c[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END c[100]
  PIN c[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END c[101]
  PIN c[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END c[102]
  PIN c[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END c[103]
  PIN c[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END c[104]
  PIN c[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END c[105]
  PIN c[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END c[106]
  PIN c[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END c[107]
  PIN c[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END c[108]
  PIN c[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END c[109]
  PIN c[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END c[10]
  PIN c[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END c[110]
  PIN c[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END c[111]
  PIN c[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END c[112]
  PIN c[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END c[113]
  PIN c[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END c[114]
  PIN c[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END c[115]
  PIN c[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END c[116]
  PIN c[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END c[117]
  PIN c[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END c[118]
  PIN c[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END c[119]
  PIN c[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END c[11]
  PIN c[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END c[120]
  PIN c[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END c[121]
  PIN c[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END c[122]
  PIN c[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END c[123]
  PIN c[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END c[124]
  PIN c[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END c[125]
  PIN c[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END c[126]
  PIN c[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END c[127]
  PIN c[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END c[12]
  PIN c[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END c[13]
  PIN c[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END c[14]
  PIN c[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END c[15]
  PIN c[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END c[16]
  PIN c[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END c[17]
  PIN c[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END c[18]
  PIN c[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END c[19]
  PIN c[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END c[1]
  PIN c[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END c[20]
  PIN c[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END c[21]
  PIN c[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END c[22]
  PIN c[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END c[23]
  PIN c[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END c[24]
  PIN c[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END c[25]
  PIN c[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END c[26]
  PIN c[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END c[27]
  PIN c[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END c[28]
  PIN c[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END c[29]
  PIN c[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END c[2]
  PIN c[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END c[30]
  PIN c[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END c[31]
  PIN c[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END c[32]
  PIN c[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END c[33]
  PIN c[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END c[34]
  PIN c[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END c[35]
  PIN c[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END c[36]
  PIN c[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END c[37]
  PIN c[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END c[38]
  PIN c[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END c[39]
  PIN c[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END c[3]
  PIN c[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END c[40]
  PIN c[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END c[41]
  PIN c[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END c[42]
  PIN c[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END c[43]
  PIN c[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END c[44]
  PIN c[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END c[45]
  PIN c[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END c[46]
  PIN c[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END c[47]
  PIN c[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END c[48]
  PIN c[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END c[49]
  PIN c[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END c[4]
  PIN c[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END c[50]
  PIN c[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END c[51]
  PIN c[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END c[52]
  PIN c[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END c[53]
  PIN c[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END c[54]
  PIN c[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END c[55]
  PIN c[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END c[56]
  PIN c[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END c[57]
  PIN c[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END c[58]
  PIN c[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END c[59]
  PIN c[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END c[5]
  PIN c[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END c[60]
  PIN c[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END c[61]
  PIN c[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END c[62]
  PIN c[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END c[63]
  PIN c[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END c[64]
  PIN c[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END c[65]
  PIN c[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END c[66]
  PIN c[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END c[67]
  PIN c[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END c[68]
  PIN c[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END c[69]
  PIN c[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END c[6]
  PIN c[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END c[70]
  PIN c[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END c[71]
  PIN c[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END c[72]
  PIN c[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END c[73]
  PIN c[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END c[74]
  PIN c[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END c[75]
  PIN c[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END c[76]
  PIN c[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END c[77]
  PIN c[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END c[78]
  PIN c[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END c[79]
  PIN c[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END c[7]
  PIN c[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END c[80]
  PIN c[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END c[81]
  PIN c[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END c[82]
  PIN c[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END c[83]
  PIN c[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END c[84]
  PIN c[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END c[85]
  PIN c[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END c[86]
  PIN c[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END c[87]
  PIN c[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END c[88]
  PIN c[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END c[89]
  PIN c[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END c[8]
  PIN c[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END c[90]
  PIN c[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END c[91]
  PIN c[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END c[92]
  PIN c[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END c[93]
  PIN c[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END c[94]
  PIN c[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END c[95]
  PIN c[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END c[96]
  PIN c[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END c[97]
  PIN c[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END c[98]
  PIN c[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END c[99]
  PIN c[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END c[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 696.000 88.440 700.000 89.040 ;
    END
  END clk
  PIN o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 696.000 26.130 700.000 ;
    END
  END o[0]
  PIN o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 531.850 696.000 532.130 700.000 ;
    END
  END o[100]
  PIN o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 536.910 696.000 537.190 700.000 ;
    END
  END o[101]
  PIN o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 541.970 696.000 542.250 700.000 ;
    END
  END o[102]
  PIN o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 547.030 696.000 547.310 700.000 ;
    END
  END o[103]
  PIN o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 552.090 696.000 552.370 700.000 ;
    END
  END o[104]
  PIN o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 557.150 696.000 557.430 700.000 ;
    END
  END o[105]
  PIN o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 562.210 696.000 562.490 700.000 ;
    END
  END o[106]
  PIN o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 567.270 696.000 567.550 700.000 ;
    END
  END o[107]
  PIN o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 572.330 696.000 572.610 700.000 ;
    END
  END o[108]
  PIN o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 577.390 696.000 577.670 700.000 ;
    END
  END o[109]
  PIN o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 696.000 76.730 700.000 ;
    END
  END o[10]
  PIN o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 582.450 696.000 582.730 700.000 ;
    END
  END o[110]
  PIN o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 587.510 696.000 587.790 700.000 ;
    END
  END o[111]
  PIN o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 592.570 696.000 592.850 700.000 ;
    END
  END o[112]
  PIN o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 597.630 696.000 597.910 700.000 ;
    END
  END o[113]
  PIN o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 602.690 696.000 602.970 700.000 ;
    END
  END o[114]
  PIN o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 607.750 696.000 608.030 700.000 ;
    END
  END o[115]
  PIN o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 612.810 696.000 613.090 700.000 ;
    END
  END o[116]
  PIN o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 617.870 696.000 618.150 700.000 ;
    END
  END o[117]
  PIN o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 622.930 696.000 623.210 700.000 ;
    END
  END o[118]
  PIN o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 627.990 696.000 628.270 700.000 ;
    END
  END o[119]
  PIN o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 696.000 81.790 700.000 ;
    END
  END o[11]
  PIN o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 633.050 696.000 633.330 700.000 ;
    END
  END o[120]
  PIN o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 638.110 696.000 638.390 700.000 ;
    END
  END o[121]
  PIN o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 643.170 696.000 643.450 700.000 ;
    END
  END o[122]
  PIN o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 648.230 696.000 648.510 700.000 ;
    END
  END o[123]
  PIN o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 653.290 696.000 653.570 700.000 ;
    END
  END o[124]
  PIN o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 658.350 696.000 658.630 700.000 ;
    END
  END o[125]
  PIN o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 663.410 696.000 663.690 700.000 ;
    END
  END o[126]
  PIN o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 668.470 696.000 668.750 700.000 ;
    END
  END o[127]
  PIN o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.570 696.000 86.850 700.000 ;
    END
  END o[12]
  PIN o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.630 696.000 91.910 700.000 ;
    END
  END o[13]
  PIN o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 696.000 96.970 700.000 ;
    END
  END o[14]
  PIN o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 696.000 102.030 700.000 ;
    END
  END o[15]
  PIN o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.810 696.000 107.090 700.000 ;
    END
  END o[16]
  PIN o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.870 696.000 112.150 700.000 ;
    END
  END o[17]
  PIN o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.930 696.000 117.210 700.000 ;
    END
  END o[18]
  PIN o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.990 696.000 122.270 700.000 ;
    END
  END o[19]
  PIN o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 30.910 696.000 31.190 700.000 ;
    END
  END o[1]
  PIN o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.050 696.000 127.330 700.000 ;
    END
  END o[20]
  PIN o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 696.000 132.390 700.000 ;
    END
  END o[21]
  PIN o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 137.170 696.000 137.450 700.000 ;
    END
  END o[22]
  PIN o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.230 696.000 142.510 700.000 ;
    END
  END o[23]
  PIN o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 696.000 147.570 700.000 ;
    END
  END o[24]
  PIN o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.350 696.000 152.630 700.000 ;
    END
  END o[25]
  PIN o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 157.410 696.000 157.690 700.000 ;
    END
  END o[26]
  PIN o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.470 696.000 162.750 700.000 ;
    END
  END o[27]
  PIN o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 696.000 167.810 700.000 ;
    END
  END o[28]
  PIN o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 172.590 696.000 172.870 700.000 ;
    END
  END o[29]
  PIN o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 696.000 36.250 700.000 ;
    END
  END o[2]
  PIN o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.650 696.000 177.930 700.000 ;
    END
  END o[30]
  PIN o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 696.000 182.990 700.000 ;
    END
  END o[31]
  PIN o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 187.770 696.000 188.050 700.000 ;
    END
  END o[32]
  PIN o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 192.830 696.000 193.110 700.000 ;
    END
  END o[33]
  PIN o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 197.890 696.000 198.170 700.000 ;
    END
  END o[34]
  PIN o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 696.000 203.230 700.000 ;
    END
  END o[35]
  PIN o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 208.010 696.000 208.290 700.000 ;
    END
  END o[36]
  PIN o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 213.070 696.000 213.350 700.000 ;
    END
  END o[37]
  PIN o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 218.130 696.000 218.410 700.000 ;
    END
  END o[38]
  PIN o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 223.190 696.000 223.470 700.000 ;
    END
  END o[39]
  PIN o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 696.000 41.310 700.000 ;
    END
  END o[3]
  PIN o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 228.250 696.000 228.530 700.000 ;
    END
  END o[40]
  PIN o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 233.310 696.000 233.590 700.000 ;
    END
  END o[41]
  PIN o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 696.000 238.650 700.000 ;
    END
  END o[42]
  PIN o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 243.430 696.000 243.710 700.000 ;
    END
  END o[43]
  PIN o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.490 696.000 248.770 700.000 ;
    END
  END o[44]
  PIN o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 253.550 696.000 253.830 700.000 ;
    END
  END o[45]
  PIN o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 258.610 696.000 258.890 700.000 ;
    END
  END o[46]
  PIN o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 263.670 696.000 263.950 700.000 ;
    END
  END o[47]
  PIN o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 268.730 696.000 269.010 700.000 ;
    END
  END o[48]
  PIN o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 273.790 696.000 274.070 700.000 ;
    END
  END o[49]
  PIN o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 696.000 46.370 700.000 ;
    END
  END o[4]
  PIN o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 278.850 696.000 279.130 700.000 ;
    END
  END o[50]
  PIN o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 283.910 696.000 284.190 700.000 ;
    END
  END o[51]
  PIN o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 288.970 696.000 289.250 700.000 ;
    END
  END o[52]
  PIN o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 294.030 696.000 294.310 700.000 ;
    END
  END o[53]
  PIN o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 299.090 696.000 299.370 700.000 ;
    END
  END o[54]
  PIN o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 304.150 696.000 304.430 700.000 ;
    END
  END o[55]
  PIN o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 309.210 696.000 309.490 700.000 ;
    END
  END o[56]
  PIN o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 314.270 696.000 314.550 700.000 ;
    END
  END o[57]
  PIN o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 319.330 696.000 319.610 700.000 ;
    END
  END o[58]
  PIN o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 324.390 696.000 324.670 700.000 ;
    END
  END o[59]
  PIN o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.150 696.000 51.430 700.000 ;
    END
  END o[5]
  PIN o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 329.450 696.000 329.730 700.000 ;
    END
  END o[60]
  PIN o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.510 696.000 334.790 700.000 ;
    END
  END o[61]
  PIN o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 339.570 696.000 339.850 700.000 ;
    END
  END o[62]
  PIN o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 696.000 344.910 700.000 ;
    END
  END o[63]
  PIN o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 349.690 696.000 349.970 700.000 ;
    END
  END o[64]
  PIN o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 354.750 696.000 355.030 700.000 ;
    END
  END o[65]
  PIN o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 359.810 696.000 360.090 700.000 ;
    END
  END o[66]
  PIN o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 364.870 696.000 365.150 700.000 ;
    END
  END o[67]
  PIN o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 369.930 696.000 370.210 700.000 ;
    END
  END o[68]
  PIN o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 374.990 696.000 375.270 700.000 ;
    END
  END o[69]
  PIN o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 696.000 56.490 700.000 ;
    END
  END o[6]
  PIN o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 380.050 696.000 380.330 700.000 ;
    END
  END o[70]
  PIN o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 385.110 696.000 385.390 700.000 ;
    END
  END o[71]
  PIN o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 390.170 696.000 390.450 700.000 ;
    END
  END o[72]
  PIN o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 395.230 696.000 395.510 700.000 ;
    END
  END o[73]
  PIN o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 400.290 696.000 400.570 700.000 ;
    END
  END o[74]
  PIN o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 405.350 696.000 405.630 700.000 ;
    END
  END o[75]
  PIN o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 410.410 696.000 410.690 700.000 ;
    END
  END o[76]
  PIN o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 415.470 696.000 415.750 700.000 ;
    END
  END o[77]
  PIN o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 420.530 696.000 420.810 700.000 ;
    END
  END o[78]
  PIN o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 425.590 696.000 425.870 700.000 ;
    END
  END o[79]
  PIN o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 696.000 61.550 700.000 ;
    END
  END o[7]
  PIN o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 430.650 696.000 430.930 700.000 ;
    END
  END o[80]
  PIN o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 435.710 696.000 435.990 700.000 ;
    END
  END o[81]
  PIN o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 440.770 696.000 441.050 700.000 ;
    END
  END o[82]
  PIN o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 445.830 696.000 446.110 700.000 ;
    END
  END o[83]
  PIN o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 450.890 696.000 451.170 700.000 ;
    END
  END o[84]
  PIN o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 455.950 696.000 456.230 700.000 ;
    END
  END o[85]
  PIN o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 461.010 696.000 461.290 700.000 ;
    END
  END o[86]
  PIN o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 466.070 696.000 466.350 700.000 ;
    END
  END o[87]
  PIN o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 471.130 696.000 471.410 700.000 ;
    END
  END o[88]
  PIN o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 476.190 696.000 476.470 700.000 ;
    END
  END o[89]
  PIN o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.330 696.000 66.610 700.000 ;
    END
  END o[8]
  PIN o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 481.250 696.000 481.530 700.000 ;
    END
  END o[90]
  PIN o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 696.000 486.590 700.000 ;
    END
  END o[91]
  PIN o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 491.370 696.000 491.650 700.000 ;
    END
  END o[92]
  PIN o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 496.430 696.000 496.710 700.000 ;
    END
  END o[93]
  PIN o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 501.490 696.000 501.770 700.000 ;
    END
  END o[94]
  PIN o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 506.550 696.000 506.830 700.000 ;
    END
  END o[95]
  PIN o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 511.610 696.000 511.890 700.000 ;
    END
  END o[96]
  PIN o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 516.670 696.000 516.950 700.000 ;
    END
  END o[97]
  PIN o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 521.730 696.000 522.010 700.000 ;
    END
  END o[98]
  PIN o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 526.790 696.000 527.070 700.000 ;
    END
  END o[99]
  PIN o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 696.000 71.670 700.000 ;
    END
  END o[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 696.000 673.810 700.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 694.330 688.350 ;
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 5.520 7.180 698.670 688.400 ;
      LAYER met2 ;
        RECT 6.080 695.720 25.570 696.730 ;
        RECT 26.410 695.720 30.630 696.730 ;
        RECT 31.470 695.720 35.690 696.730 ;
        RECT 36.530 695.720 40.750 696.730 ;
        RECT 41.590 695.720 45.810 696.730 ;
        RECT 46.650 695.720 50.870 696.730 ;
        RECT 51.710 695.720 55.930 696.730 ;
        RECT 56.770 695.720 60.990 696.730 ;
        RECT 61.830 695.720 66.050 696.730 ;
        RECT 66.890 695.720 71.110 696.730 ;
        RECT 71.950 695.720 76.170 696.730 ;
        RECT 77.010 695.720 81.230 696.730 ;
        RECT 82.070 695.720 86.290 696.730 ;
        RECT 87.130 695.720 91.350 696.730 ;
        RECT 92.190 695.720 96.410 696.730 ;
        RECT 97.250 695.720 101.470 696.730 ;
        RECT 102.310 695.720 106.530 696.730 ;
        RECT 107.370 695.720 111.590 696.730 ;
        RECT 112.430 695.720 116.650 696.730 ;
        RECT 117.490 695.720 121.710 696.730 ;
        RECT 122.550 695.720 126.770 696.730 ;
        RECT 127.610 695.720 131.830 696.730 ;
        RECT 132.670 695.720 136.890 696.730 ;
        RECT 137.730 695.720 141.950 696.730 ;
        RECT 142.790 695.720 147.010 696.730 ;
        RECT 147.850 695.720 152.070 696.730 ;
        RECT 152.910 695.720 157.130 696.730 ;
        RECT 157.970 695.720 162.190 696.730 ;
        RECT 163.030 695.720 167.250 696.730 ;
        RECT 168.090 695.720 172.310 696.730 ;
        RECT 173.150 695.720 177.370 696.730 ;
        RECT 178.210 695.720 182.430 696.730 ;
        RECT 183.270 695.720 187.490 696.730 ;
        RECT 188.330 695.720 192.550 696.730 ;
        RECT 193.390 695.720 197.610 696.730 ;
        RECT 198.450 695.720 202.670 696.730 ;
        RECT 203.510 695.720 207.730 696.730 ;
        RECT 208.570 695.720 212.790 696.730 ;
        RECT 213.630 695.720 217.850 696.730 ;
        RECT 218.690 695.720 222.910 696.730 ;
        RECT 223.750 695.720 227.970 696.730 ;
        RECT 228.810 695.720 233.030 696.730 ;
        RECT 233.870 695.720 238.090 696.730 ;
        RECT 238.930 695.720 243.150 696.730 ;
        RECT 243.990 695.720 248.210 696.730 ;
        RECT 249.050 695.720 253.270 696.730 ;
        RECT 254.110 695.720 258.330 696.730 ;
        RECT 259.170 695.720 263.390 696.730 ;
        RECT 264.230 695.720 268.450 696.730 ;
        RECT 269.290 695.720 273.510 696.730 ;
        RECT 274.350 695.720 278.570 696.730 ;
        RECT 279.410 695.720 283.630 696.730 ;
        RECT 284.470 695.720 288.690 696.730 ;
        RECT 289.530 695.720 293.750 696.730 ;
        RECT 294.590 695.720 298.810 696.730 ;
        RECT 299.650 695.720 303.870 696.730 ;
        RECT 304.710 695.720 308.930 696.730 ;
        RECT 309.770 695.720 313.990 696.730 ;
        RECT 314.830 695.720 319.050 696.730 ;
        RECT 319.890 695.720 324.110 696.730 ;
        RECT 324.950 695.720 329.170 696.730 ;
        RECT 330.010 695.720 334.230 696.730 ;
        RECT 335.070 695.720 339.290 696.730 ;
        RECT 340.130 695.720 344.350 696.730 ;
        RECT 345.190 695.720 349.410 696.730 ;
        RECT 350.250 695.720 354.470 696.730 ;
        RECT 355.310 695.720 359.530 696.730 ;
        RECT 360.370 695.720 364.590 696.730 ;
        RECT 365.430 695.720 369.650 696.730 ;
        RECT 370.490 695.720 374.710 696.730 ;
        RECT 375.550 695.720 379.770 696.730 ;
        RECT 380.610 695.720 384.830 696.730 ;
        RECT 385.670 695.720 389.890 696.730 ;
        RECT 390.730 695.720 394.950 696.730 ;
        RECT 395.790 695.720 400.010 696.730 ;
        RECT 400.850 695.720 405.070 696.730 ;
        RECT 405.910 695.720 410.130 696.730 ;
        RECT 410.970 695.720 415.190 696.730 ;
        RECT 416.030 695.720 420.250 696.730 ;
        RECT 421.090 695.720 425.310 696.730 ;
        RECT 426.150 695.720 430.370 696.730 ;
        RECT 431.210 695.720 435.430 696.730 ;
        RECT 436.270 695.720 440.490 696.730 ;
        RECT 441.330 695.720 445.550 696.730 ;
        RECT 446.390 695.720 450.610 696.730 ;
        RECT 451.450 695.720 455.670 696.730 ;
        RECT 456.510 695.720 460.730 696.730 ;
        RECT 461.570 695.720 465.790 696.730 ;
        RECT 466.630 695.720 470.850 696.730 ;
        RECT 471.690 695.720 475.910 696.730 ;
        RECT 476.750 695.720 480.970 696.730 ;
        RECT 481.810 695.720 486.030 696.730 ;
        RECT 486.870 695.720 491.090 696.730 ;
        RECT 491.930 695.720 496.150 696.730 ;
        RECT 496.990 695.720 501.210 696.730 ;
        RECT 502.050 695.720 506.270 696.730 ;
        RECT 507.110 695.720 511.330 696.730 ;
        RECT 512.170 695.720 516.390 696.730 ;
        RECT 517.230 695.720 521.450 696.730 ;
        RECT 522.290 695.720 526.510 696.730 ;
        RECT 527.350 695.720 531.570 696.730 ;
        RECT 532.410 695.720 536.630 696.730 ;
        RECT 537.470 695.720 541.690 696.730 ;
        RECT 542.530 695.720 546.750 696.730 ;
        RECT 547.590 695.720 551.810 696.730 ;
        RECT 552.650 695.720 556.870 696.730 ;
        RECT 557.710 695.720 561.930 696.730 ;
        RECT 562.770 695.720 566.990 696.730 ;
        RECT 567.830 695.720 572.050 696.730 ;
        RECT 572.890 695.720 577.110 696.730 ;
        RECT 577.950 695.720 582.170 696.730 ;
        RECT 583.010 695.720 587.230 696.730 ;
        RECT 588.070 695.720 592.290 696.730 ;
        RECT 593.130 695.720 597.350 696.730 ;
        RECT 598.190 695.720 602.410 696.730 ;
        RECT 603.250 695.720 607.470 696.730 ;
        RECT 608.310 695.720 612.530 696.730 ;
        RECT 613.370 695.720 617.590 696.730 ;
        RECT 618.430 695.720 622.650 696.730 ;
        RECT 623.490 695.720 627.710 696.730 ;
        RECT 628.550 695.720 632.770 696.730 ;
        RECT 633.610 695.720 637.830 696.730 ;
        RECT 638.670 695.720 642.890 696.730 ;
        RECT 643.730 695.720 647.950 696.730 ;
        RECT 648.790 695.720 653.010 696.730 ;
        RECT 653.850 695.720 658.070 696.730 ;
        RECT 658.910 695.720 663.130 696.730 ;
        RECT 663.970 695.720 668.190 696.730 ;
        RECT 669.030 695.720 673.250 696.730 ;
        RECT 674.090 695.720 698.650 696.730 ;
        RECT 6.080 4.280 698.650 695.720 ;
        RECT 6.080 3.670 28.330 4.280 ;
        RECT 29.170 3.670 33.390 4.280 ;
        RECT 34.230 3.670 38.450 4.280 ;
        RECT 39.290 3.670 43.510 4.280 ;
        RECT 44.350 3.670 48.570 4.280 ;
        RECT 49.410 3.670 53.630 4.280 ;
        RECT 54.470 3.670 58.690 4.280 ;
        RECT 59.530 3.670 63.750 4.280 ;
        RECT 64.590 3.670 68.810 4.280 ;
        RECT 69.650 3.670 73.870 4.280 ;
        RECT 74.710 3.670 78.930 4.280 ;
        RECT 79.770 3.670 83.990 4.280 ;
        RECT 84.830 3.670 89.050 4.280 ;
        RECT 89.890 3.670 94.110 4.280 ;
        RECT 94.950 3.670 99.170 4.280 ;
        RECT 100.010 3.670 104.230 4.280 ;
        RECT 105.070 3.670 109.290 4.280 ;
        RECT 110.130 3.670 114.350 4.280 ;
        RECT 115.190 3.670 119.410 4.280 ;
        RECT 120.250 3.670 124.470 4.280 ;
        RECT 125.310 3.670 129.530 4.280 ;
        RECT 130.370 3.670 134.590 4.280 ;
        RECT 135.430 3.670 139.650 4.280 ;
        RECT 140.490 3.670 144.710 4.280 ;
        RECT 145.550 3.670 149.770 4.280 ;
        RECT 150.610 3.670 154.830 4.280 ;
        RECT 155.670 3.670 159.890 4.280 ;
        RECT 160.730 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.010 4.280 ;
        RECT 170.850 3.670 175.070 4.280 ;
        RECT 175.910 3.670 180.130 4.280 ;
        RECT 180.970 3.670 185.190 4.280 ;
        RECT 186.030 3.670 190.250 4.280 ;
        RECT 191.090 3.670 195.310 4.280 ;
        RECT 196.150 3.670 200.370 4.280 ;
        RECT 201.210 3.670 205.430 4.280 ;
        RECT 206.270 3.670 210.490 4.280 ;
        RECT 211.330 3.670 215.550 4.280 ;
        RECT 216.390 3.670 220.610 4.280 ;
        RECT 221.450 3.670 225.670 4.280 ;
        RECT 226.510 3.670 230.730 4.280 ;
        RECT 231.570 3.670 235.790 4.280 ;
        RECT 236.630 3.670 240.850 4.280 ;
        RECT 241.690 3.670 245.910 4.280 ;
        RECT 246.750 3.670 250.970 4.280 ;
        RECT 251.810 3.670 256.030 4.280 ;
        RECT 256.870 3.670 261.090 4.280 ;
        RECT 261.930 3.670 266.150 4.280 ;
        RECT 266.990 3.670 271.210 4.280 ;
        RECT 272.050 3.670 276.270 4.280 ;
        RECT 277.110 3.670 281.330 4.280 ;
        RECT 282.170 3.670 286.390 4.280 ;
        RECT 287.230 3.670 291.450 4.280 ;
        RECT 292.290 3.670 296.510 4.280 ;
        RECT 297.350 3.670 301.570 4.280 ;
        RECT 302.410 3.670 306.630 4.280 ;
        RECT 307.470 3.670 311.690 4.280 ;
        RECT 312.530 3.670 316.750 4.280 ;
        RECT 317.590 3.670 321.810 4.280 ;
        RECT 322.650 3.670 326.870 4.280 ;
        RECT 327.710 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.990 4.280 ;
        RECT 337.830 3.670 342.050 4.280 ;
        RECT 342.890 3.670 347.110 4.280 ;
        RECT 347.950 3.670 352.170 4.280 ;
        RECT 353.010 3.670 357.230 4.280 ;
        RECT 358.070 3.670 362.290 4.280 ;
        RECT 363.130 3.670 367.350 4.280 ;
        RECT 368.190 3.670 372.410 4.280 ;
        RECT 373.250 3.670 377.470 4.280 ;
        RECT 378.310 3.670 382.530 4.280 ;
        RECT 383.370 3.670 387.590 4.280 ;
        RECT 388.430 3.670 392.650 4.280 ;
        RECT 393.490 3.670 397.710 4.280 ;
        RECT 398.550 3.670 402.770 4.280 ;
        RECT 403.610 3.670 407.830 4.280 ;
        RECT 408.670 3.670 412.890 4.280 ;
        RECT 413.730 3.670 417.950 4.280 ;
        RECT 418.790 3.670 423.010 4.280 ;
        RECT 423.850 3.670 428.070 4.280 ;
        RECT 428.910 3.670 433.130 4.280 ;
        RECT 433.970 3.670 438.190 4.280 ;
        RECT 439.030 3.670 443.250 4.280 ;
        RECT 444.090 3.670 448.310 4.280 ;
        RECT 449.150 3.670 453.370 4.280 ;
        RECT 454.210 3.670 458.430 4.280 ;
        RECT 459.270 3.670 463.490 4.280 ;
        RECT 464.330 3.670 468.550 4.280 ;
        RECT 469.390 3.670 473.610 4.280 ;
        RECT 474.450 3.670 478.670 4.280 ;
        RECT 479.510 3.670 483.730 4.280 ;
        RECT 484.570 3.670 488.790 4.280 ;
        RECT 489.630 3.670 493.850 4.280 ;
        RECT 494.690 3.670 498.910 4.280 ;
        RECT 499.750 3.670 503.970 4.280 ;
        RECT 504.810 3.670 509.030 4.280 ;
        RECT 509.870 3.670 514.090 4.280 ;
        RECT 514.930 3.670 519.150 4.280 ;
        RECT 519.990 3.670 524.210 4.280 ;
        RECT 525.050 3.670 529.270 4.280 ;
        RECT 530.110 3.670 534.330 4.280 ;
        RECT 535.170 3.670 539.390 4.280 ;
        RECT 540.230 3.670 544.450 4.280 ;
        RECT 545.290 3.670 549.510 4.280 ;
        RECT 550.350 3.670 554.570 4.280 ;
        RECT 555.410 3.670 559.630 4.280 ;
        RECT 560.470 3.670 564.690 4.280 ;
        RECT 565.530 3.670 569.750 4.280 ;
        RECT 570.590 3.670 574.810 4.280 ;
        RECT 575.650 3.670 579.870 4.280 ;
        RECT 580.710 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.990 4.280 ;
        RECT 590.830 3.670 595.050 4.280 ;
        RECT 595.890 3.670 600.110 4.280 ;
        RECT 600.950 3.670 605.170 4.280 ;
        RECT 606.010 3.670 610.230 4.280 ;
        RECT 611.070 3.670 615.290 4.280 ;
        RECT 616.130 3.670 620.350 4.280 ;
        RECT 621.190 3.670 625.410 4.280 ;
        RECT 626.250 3.670 630.470 4.280 ;
        RECT 631.310 3.670 635.530 4.280 ;
        RECT 636.370 3.670 640.590 4.280 ;
        RECT 641.430 3.670 645.650 4.280 ;
        RECT 646.490 3.670 650.710 4.280 ;
        RECT 651.550 3.670 655.770 4.280 ;
        RECT 656.610 3.670 660.830 4.280 ;
        RECT 661.670 3.670 665.890 4.280 ;
        RECT 666.730 3.670 670.950 4.280 ;
        RECT 671.790 3.670 698.650 4.280 ;
      LAYER met3 ;
        RECT 9.130 611.680 698.675 688.325 ;
        RECT 9.130 610.280 695.600 611.680 ;
        RECT 9.130 607.600 698.675 610.280 ;
        RECT 9.130 606.200 695.600 607.600 ;
        RECT 9.130 603.520 698.675 606.200 ;
        RECT 9.130 602.120 695.600 603.520 ;
        RECT 9.130 599.440 698.675 602.120 ;
        RECT 9.130 598.040 695.600 599.440 ;
        RECT 9.130 595.360 698.675 598.040 ;
        RECT 9.130 593.960 695.600 595.360 ;
        RECT 9.130 591.280 698.675 593.960 ;
        RECT 9.130 589.880 695.600 591.280 ;
        RECT 9.130 587.200 698.675 589.880 ;
        RECT 9.130 585.800 695.600 587.200 ;
        RECT 9.130 583.120 698.675 585.800 ;
        RECT 9.130 581.720 695.600 583.120 ;
        RECT 9.130 579.040 698.675 581.720 ;
        RECT 9.130 577.640 695.600 579.040 ;
        RECT 9.130 574.960 698.675 577.640 ;
        RECT 9.130 573.560 695.600 574.960 ;
        RECT 9.130 570.880 698.675 573.560 ;
        RECT 9.130 569.480 695.600 570.880 ;
        RECT 9.130 566.800 698.675 569.480 ;
        RECT 9.130 565.400 695.600 566.800 ;
        RECT 9.130 562.720 698.675 565.400 ;
        RECT 9.130 561.320 695.600 562.720 ;
        RECT 9.130 558.640 698.675 561.320 ;
        RECT 9.130 557.240 695.600 558.640 ;
        RECT 9.130 554.560 698.675 557.240 ;
        RECT 9.130 553.160 695.600 554.560 ;
        RECT 9.130 550.480 698.675 553.160 ;
        RECT 9.130 549.080 695.600 550.480 ;
        RECT 9.130 546.400 698.675 549.080 ;
        RECT 9.130 545.000 695.600 546.400 ;
        RECT 9.130 542.320 698.675 545.000 ;
        RECT 9.130 540.920 695.600 542.320 ;
        RECT 9.130 538.240 698.675 540.920 ;
        RECT 9.130 536.840 695.600 538.240 ;
        RECT 9.130 534.160 698.675 536.840 ;
        RECT 9.130 532.760 695.600 534.160 ;
        RECT 9.130 530.080 698.675 532.760 ;
        RECT 9.130 528.680 695.600 530.080 ;
        RECT 9.130 526.000 698.675 528.680 ;
        RECT 9.130 524.600 695.600 526.000 ;
        RECT 9.130 521.920 698.675 524.600 ;
        RECT 9.130 520.520 695.600 521.920 ;
        RECT 9.130 517.840 698.675 520.520 ;
        RECT 9.130 516.440 695.600 517.840 ;
        RECT 9.130 513.760 698.675 516.440 ;
        RECT 9.130 512.360 695.600 513.760 ;
        RECT 9.130 509.680 698.675 512.360 ;
        RECT 9.130 508.280 695.600 509.680 ;
        RECT 9.130 505.600 698.675 508.280 ;
        RECT 9.130 504.200 695.600 505.600 ;
        RECT 9.130 501.520 698.675 504.200 ;
        RECT 9.130 500.120 695.600 501.520 ;
        RECT 9.130 497.440 698.675 500.120 ;
        RECT 9.130 496.040 695.600 497.440 ;
        RECT 9.130 493.360 698.675 496.040 ;
        RECT 9.130 491.960 695.600 493.360 ;
        RECT 9.130 489.280 698.675 491.960 ;
        RECT 9.130 487.880 695.600 489.280 ;
        RECT 9.130 485.200 698.675 487.880 ;
        RECT 9.130 483.800 695.600 485.200 ;
        RECT 9.130 481.120 698.675 483.800 ;
        RECT 9.130 479.720 695.600 481.120 ;
        RECT 9.130 477.040 698.675 479.720 ;
        RECT 9.130 475.640 695.600 477.040 ;
        RECT 9.130 472.960 698.675 475.640 ;
        RECT 9.130 471.560 695.600 472.960 ;
        RECT 9.130 468.880 698.675 471.560 ;
        RECT 9.130 467.480 695.600 468.880 ;
        RECT 9.130 464.800 698.675 467.480 ;
        RECT 9.130 463.400 695.600 464.800 ;
        RECT 9.130 460.720 698.675 463.400 ;
        RECT 9.130 459.320 695.600 460.720 ;
        RECT 9.130 456.640 698.675 459.320 ;
        RECT 9.130 455.240 695.600 456.640 ;
        RECT 9.130 452.560 698.675 455.240 ;
        RECT 9.130 451.160 695.600 452.560 ;
        RECT 9.130 448.480 698.675 451.160 ;
        RECT 9.130 447.080 695.600 448.480 ;
        RECT 9.130 444.400 698.675 447.080 ;
        RECT 9.130 443.000 695.600 444.400 ;
        RECT 9.130 440.320 698.675 443.000 ;
        RECT 9.130 438.920 695.600 440.320 ;
        RECT 9.130 436.240 698.675 438.920 ;
        RECT 9.130 434.840 695.600 436.240 ;
        RECT 9.130 432.160 698.675 434.840 ;
        RECT 9.130 430.760 695.600 432.160 ;
        RECT 9.130 428.080 698.675 430.760 ;
        RECT 9.130 426.680 695.600 428.080 ;
        RECT 9.130 424.000 698.675 426.680 ;
        RECT 9.130 422.600 695.600 424.000 ;
        RECT 9.130 419.920 698.675 422.600 ;
        RECT 9.130 418.520 695.600 419.920 ;
        RECT 9.130 415.840 698.675 418.520 ;
        RECT 9.130 414.440 695.600 415.840 ;
        RECT 9.130 411.760 698.675 414.440 ;
        RECT 9.130 410.360 695.600 411.760 ;
        RECT 9.130 407.680 698.675 410.360 ;
        RECT 9.130 406.280 695.600 407.680 ;
        RECT 9.130 403.600 698.675 406.280 ;
        RECT 9.130 402.200 695.600 403.600 ;
        RECT 9.130 399.520 698.675 402.200 ;
        RECT 9.130 398.120 695.600 399.520 ;
        RECT 9.130 395.440 698.675 398.120 ;
        RECT 9.130 394.040 695.600 395.440 ;
        RECT 9.130 391.360 698.675 394.040 ;
        RECT 9.130 389.960 695.600 391.360 ;
        RECT 9.130 387.280 698.675 389.960 ;
        RECT 9.130 385.880 695.600 387.280 ;
        RECT 9.130 383.200 698.675 385.880 ;
        RECT 9.130 381.800 695.600 383.200 ;
        RECT 9.130 379.120 698.675 381.800 ;
        RECT 9.130 377.720 695.600 379.120 ;
        RECT 9.130 375.040 698.675 377.720 ;
        RECT 9.130 373.640 695.600 375.040 ;
        RECT 9.130 370.960 698.675 373.640 ;
        RECT 9.130 369.560 695.600 370.960 ;
        RECT 9.130 366.880 698.675 369.560 ;
        RECT 9.130 365.480 695.600 366.880 ;
        RECT 9.130 362.800 698.675 365.480 ;
        RECT 9.130 361.400 695.600 362.800 ;
        RECT 9.130 358.720 698.675 361.400 ;
        RECT 9.130 357.320 695.600 358.720 ;
        RECT 9.130 354.640 698.675 357.320 ;
        RECT 9.130 353.240 695.600 354.640 ;
        RECT 9.130 350.560 698.675 353.240 ;
        RECT 9.130 349.160 695.600 350.560 ;
        RECT 9.130 346.480 698.675 349.160 ;
        RECT 9.130 345.080 695.600 346.480 ;
        RECT 9.130 342.400 698.675 345.080 ;
        RECT 9.130 341.000 695.600 342.400 ;
        RECT 9.130 338.320 698.675 341.000 ;
        RECT 9.130 336.920 695.600 338.320 ;
        RECT 9.130 334.240 698.675 336.920 ;
        RECT 9.130 332.840 695.600 334.240 ;
        RECT 9.130 330.160 698.675 332.840 ;
        RECT 9.130 328.760 695.600 330.160 ;
        RECT 9.130 326.080 698.675 328.760 ;
        RECT 9.130 324.680 695.600 326.080 ;
        RECT 9.130 322.000 698.675 324.680 ;
        RECT 9.130 320.600 695.600 322.000 ;
        RECT 9.130 317.920 698.675 320.600 ;
        RECT 9.130 316.520 695.600 317.920 ;
        RECT 9.130 313.840 698.675 316.520 ;
        RECT 9.130 312.440 695.600 313.840 ;
        RECT 9.130 309.760 698.675 312.440 ;
        RECT 9.130 308.360 695.600 309.760 ;
        RECT 9.130 305.680 698.675 308.360 ;
        RECT 9.130 304.280 695.600 305.680 ;
        RECT 9.130 301.600 698.675 304.280 ;
        RECT 9.130 300.200 695.600 301.600 ;
        RECT 9.130 297.520 698.675 300.200 ;
        RECT 9.130 296.120 695.600 297.520 ;
        RECT 9.130 293.440 698.675 296.120 ;
        RECT 9.130 292.040 695.600 293.440 ;
        RECT 9.130 289.360 698.675 292.040 ;
        RECT 9.130 287.960 695.600 289.360 ;
        RECT 9.130 285.280 698.675 287.960 ;
        RECT 9.130 283.880 695.600 285.280 ;
        RECT 9.130 281.200 698.675 283.880 ;
        RECT 9.130 279.800 695.600 281.200 ;
        RECT 9.130 277.120 698.675 279.800 ;
        RECT 9.130 275.720 695.600 277.120 ;
        RECT 9.130 273.040 698.675 275.720 ;
        RECT 9.130 271.640 695.600 273.040 ;
        RECT 9.130 268.960 698.675 271.640 ;
        RECT 9.130 267.560 695.600 268.960 ;
        RECT 9.130 264.880 698.675 267.560 ;
        RECT 9.130 263.480 695.600 264.880 ;
        RECT 9.130 260.800 698.675 263.480 ;
        RECT 9.130 259.400 695.600 260.800 ;
        RECT 9.130 256.720 698.675 259.400 ;
        RECT 9.130 255.320 695.600 256.720 ;
        RECT 9.130 252.640 698.675 255.320 ;
        RECT 9.130 251.240 695.600 252.640 ;
        RECT 9.130 248.560 698.675 251.240 ;
        RECT 9.130 247.160 695.600 248.560 ;
        RECT 9.130 244.480 698.675 247.160 ;
        RECT 9.130 243.080 695.600 244.480 ;
        RECT 9.130 240.400 698.675 243.080 ;
        RECT 9.130 239.000 695.600 240.400 ;
        RECT 9.130 236.320 698.675 239.000 ;
        RECT 9.130 234.920 695.600 236.320 ;
        RECT 9.130 232.240 698.675 234.920 ;
        RECT 9.130 230.840 695.600 232.240 ;
        RECT 9.130 228.160 698.675 230.840 ;
        RECT 9.130 226.760 695.600 228.160 ;
        RECT 9.130 224.080 698.675 226.760 ;
        RECT 9.130 222.680 695.600 224.080 ;
        RECT 9.130 220.000 698.675 222.680 ;
        RECT 9.130 218.600 695.600 220.000 ;
        RECT 9.130 215.920 698.675 218.600 ;
        RECT 9.130 214.520 695.600 215.920 ;
        RECT 9.130 211.840 698.675 214.520 ;
        RECT 9.130 210.440 695.600 211.840 ;
        RECT 9.130 207.760 698.675 210.440 ;
        RECT 9.130 206.360 695.600 207.760 ;
        RECT 9.130 203.680 698.675 206.360 ;
        RECT 9.130 202.280 695.600 203.680 ;
        RECT 9.130 199.600 698.675 202.280 ;
        RECT 9.130 198.200 695.600 199.600 ;
        RECT 9.130 195.520 698.675 198.200 ;
        RECT 9.130 194.120 695.600 195.520 ;
        RECT 9.130 191.440 698.675 194.120 ;
        RECT 9.130 190.040 695.600 191.440 ;
        RECT 9.130 187.360 698.675 190.040 ;
        RECT 9.130 185.960 695.600 187.360 ;
        RECT 9.130 183.280 698.675 185.960 ;
        RECT 9.130 181.880 695.600 183.280 ;
        RECT 9.130 179.200 698.675 181.880 ;
        RECT 9.130 177.800 695.600 179.200 ;
        RECT 9.130 175.120 698.675 177.800 ;
        RECT 9.130 173.720 695.600 175.120 ;
        RECT 9.130 171.040 698.675 173.720 ;
        RECT 9.130 169.640 695.600 171.040 ;
        RECT 9.130 166.960 698.675 169.640 ;
        RECT 9.130 165.560 695.600 166.960 ;
        RECT 9.130 162.880 698.675 165.560 ;
        RECT 9.130 161.480 695.600 162.880 ;
        RECT 9.130 158.800 698.675 161.480 ;
        RECT 9.130 157.400 695.600 158.800 ;
        RECT 9.130 154.720 698.675 157.400 ;
        RECT 9.130 153.320 695.600 154.720 ;
        RECT 9.130 150.640 698.675 153.320 ;
        RECT 9.130 149.240 695.600 150.640 ;
        RECT 9.130 146.560 698.675 149.240 ;
        RECT 9.130 145.160 695.600 146.560 ;
        RECT 9.130 142.480 698.675 145.160 ;
        RECT 9.130 141.080 695.600 142.480 ;
        RECT 9.130 138.400 698.675 141.080 ;
        RECT 9.130 137.000 695.600 138.400 ;
        RECT 9.130 134.320 698.675 137.000 ;
        RECT 9.130 132.920 695.600 134.320 ;
        RECT 9.130 130.240 698.675 132.920 ;
        RECT 9.130 128.840 695.600 130.240 ;
        RECT 9.130 126.160 698.675 128.840 ;
        RECT 9.130 124.760 695.600 126.160 ;
        RECT 9.130 122.080 698.675 124.760 ;
        RECT 9.130 120.680 695.600 122.080 ;
        RECT 9.130 118.000 698.675 120.680 ;
        RECT 9.130 116.600 695.600 118.000 ;
        RECT 9.130 113.920 698.675 116.600 ;
        RECT 9.130 112.520 695.600 113.920 ;
        RECT 9.130 109.840 698.675 112.520 ;
        RECT 9.130 108.440 695.600 109.840 ;
        RECT 9.130 105.760 698.675 108.440 ;
        RECT 9.130 104.360 695.600 105.760 ;
        RECT 9.130 101.680 698.675 104.360 ;
        RECT 9.130 100.280 695.600 101.680 ;
        RECT 9.130 97.600 698.675 100.280 ;
        RECT 9.130 96.200 695.600 97.600 ;
        RECT 9.130 93.520 698.675 96.200 ;
        RECT 9.130 92.120 695.600 93.520 ;
        RECT 9.130 89.440 698.675 92.120 ;
        RECT 9.130 88.040 695.600 89.440 ;
        RECT 9.130 10.715 698.675 88.040 ;
      LAYER met4 ;
        RECT 19.615 13.775 27.170 669.625 ;
        RECT 31.070 13.775 188.570 669.625 ;
        RECT 192.470 13.775 207.170 669.625 ;
        RECT 211.070 13.775 368.570 669.625 ;
        RECT 372.470 13.775 387.170 669.625 ;
        RECT 391.070 13.775 548.570 669.625 ;
        RECT 552.470 13.775 567.170 669.625 ;
        RECT 571.070 13.775 690.625 669.625 ;
  END
END multiply_add_64x64
END LIBRARY

