* NGSPICE file created from Microwatt_FP_DFFRFile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

.subckt Microwatt_FP_DFFRFile CLK D1[0] D1[10] D1[11] D1[12] D1[13] D1[14] D1[15]
+ D1[16] D1[17] D1[18] D1[19] D1[1] D1[20] D1[21] D1[22] D1[23] D1[24] D1[25] D1[26]
+ D1[27] D1[28] D1[29] D1[2] D1[30] D1[31] D1[32] D1[33] D1[34] D1[35] D1[36] D1[37]
+ D1[38] D1[39] D1[3] D1[40] D1[41] D1[42] D1[43] D1[44] D1[45] D1[46] D1[47] D1[48]
+ D1[49] D1[4] D1[50] D1[51] D1[52] D1[53] D1[54] D1[55] D1[56] D1[57] D1[58] D1[59]
+ D1[5] D1[60] D1[61] D1[62] D1[63] D1[6] D1[7] D1[8] D1[9] D2[0] D2[10] D2[11] D2[12]
+ D2[13] D2[14] D2[15] D2[16] D2[17] D2[18] D2[19] D2[1] D2[20] D2[21] D2[22] D2[23]
+ D2[24] D2[25] D2[26] D2[27] D2[28] D2[29] D2[2] D2[30] D2[31] D2[32] D2[33] D2[34]
+ D2[35] D2[36] D2[37] D2[38] D2[39] D2[3] D2[40] D2[41] D2[42] D2[43] D2[44] D2[45]
+ D2[46] D2[47] D2[48] D2[49] D2[4] D2[50] D2[51] D2[52] D2[53] D2[54] D2[55] D2[56]
+ D2[57] D2[58] D2[59] D2[5] D2[60] D2[61] D2[62] D2[63] D2[6] D2[7] D2[8] D2[9] D3[0]
+ D3[10] D3[11] D3[12] D3[13] D3[14] D3[15] D3[16] D3[17] D3[18] D3[19] D3[1] D3[20]
+ D3[21] D3[22] D3[23] D3[24] D3[25] D3[26] D3[27] D3[28] D3[29] D3[2] D3[30] D3[31]
+ D3[32] D3[33] D3[34] D3[35] D3[36] D3[37] D3[38] D3[39] D3[3] D3[40] D3[41] D3[42]
+ D3[43] D3[44] D3[45] D3[46] D3[47] D3[48] D3[49] D3[4] D3[50] D3[51] D3[52] D3[53]
+ D3[54] D3[55] D3[56] D3[57] D3[58] D3[59] D3[5] D3[60] D3[61] D3[62] D3[63] D3[6]
+ D3[7] D3[8] D3[9] DW[0] DW[10] DW[11] DW[12] DW[13] DW[14] DW[15] DW[16] DW[17]
+ DW[18] DW[19] DW[1] DW[20] DW[21] DW[22] DW[23] DW[24] DW[25] DW[26] DW[27] DW[28]
+ DW[29] DW[2] DW[30] DW[31] DW[32] DW[33] DW[34] DW[35] DW[36] DW[37] DW[38] DW[39]
+ DW[3] DW[40] DW[41] DW[42] DW[43] DW[44] DW[45] DW[46] DW[47] DW[48] DW[49] DW[4]
+ DW[50] DW[51] DW[52] DW[53] DW[54] DW[55] DW[56] DW[57] DW[58] DW[59] DW[5] DW[60]
+ DW[61] DW[62] DW[63] DW[6] DW[7] DW[8] DW[9] R1[0] R1[1] R1[2] R1[3] R1[4] R1[5]
+ R2[0] R2[1] R2[2] R2[3] R2[4] R2[5] R3[0] R3[1] R3[2] R3[3] R3[4] R3[5] RW[0] RW[1]
+ RW[2] RW[3] RW[4] RW[5] VGND VPWR WE
XFILLER_228_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34984_ clknet_leaf_457_CLK _03098_ VGND VGND VPWR VPWR registers\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1360 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1371 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1382 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33935_ clknet_leaf_133_CLK _02049_ VGND VGND VPWR VPWR registers\[37\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1393 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18869_ _05404_ _05616_ _05617_ _05410_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__a22o_1
XFILLER_55_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20900_ _07377_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__buf_6
X_21880_ _08540_ _08544_ _08405_ _08406_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__o211a_1
X_33866_ clknet_leaf_153_CLK _01980_ VGND VGND VPWR VPWR registers\[3\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35605_ clknet_leaf_79_CLK _03719_ VGND VGND VPWR VPWR registers\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_20831_ registers\[24\]\[4\] registers\[25\]\[4\] registers\[26\]\[4\] registers\[27\]\[4\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__mux4_1
X_32817_ clknet_leaf_367_CLK _00931_ VGND VGND VPWR VPWR registers\[55\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33797_ clknet_leaf_250_CLK _01911_ VGND VGND VPWR VPWR registers\[40\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23550_ _09934_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__clkbuf_1
X_35536_ clknet_leaf_138_CLK _03650_ VGND VGND VPWR VPWR registers\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_20762_ _07455_ _07458_ _07370_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__o21ba_1
X_32748_ clknet_leaf_371_CLK _00862_ VGND VGND VPWR VPWR registers\[56\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_22501_ _07312_ VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__buf_4
XFILLER_126_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23481_ _09898_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
X_35467_ clknet_leaf_150_CLK _03581_ VGND VGND VPWR VPWR registers\[14\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20693_ _07328_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__buf_12
XFILLER_56_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32679_ clknet_leaf_436_CLK _00793_ VGND VGND VPWR VPWR registers\[57\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22432_ registers\[36\]\[50\] registers\[37\]\[50\] registers\[38\]\[50\] registers\[39\]\[50\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__mux4_1
X_25220_ _10760_ registers\[51\]\[14\] _10876_ VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34418_ clknet_leaf_411_CLK _02532_ VGND VGND VPWR VPWR registers\[30\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35398_ clknet_leaf_215_CLK _03512_ VGND VGND VPWR VPWR registers\[15\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25151_ _10838_ registers\[52\]\[51\] _10836_ VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__mux2_1
X_22363_ registers\[56\]\[48\] registers\[57\]\[48\] registers\[58\]\[48\] registers\[59\]\[48\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__mux4_1
XFILLER_52_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34349_ clknet_leaf_403_CLK _02463_ VGND VGND VPWR VPWR registers\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_248_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24102_ _09642_ registers\[5\]\[61\] _10160_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__mux2_1
X_21314_ _07301_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25082_ _10791_ registers\[52\]\[29\] _10773_ VGND VGND VPWR VPWR _10792_ sky130_fd_sc_hd__mux2_1
XFILLER_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22294_ registers\[60\]\[46\] registers\[61\]\[46\] registers\[62\]\[46\] registers\[63\]\[46\]
+ _08884_ _08678_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__mux4_1
X_28910_ _12858_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__clkbuf_1
X_24033_ _09573_ registers\[5\]\[28\] _10183_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__mux2_1
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21245_ _07924_ _07925_ _07926_ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__a22o_1
X_36019_ clknet_leaf_356_CLK _04133_ VGND VGND VPWR VPWR registers\[63\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29890_ _13405_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28841_ _12822_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21176_ registers\[0\]\[14\] registers\[1\]\[14\] registers\[2\]\[14\] registers\[3\]\[14\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__mux4_1
XFILLER_81_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20127_ registers\[32\]\[50\] registers\[33\]\[50\] registers\[34\]\[50\] registers\[35\]\[50\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28772_ _11857_ registers\[26\]\[61\] _12718_ VGND VGND VPWR VPWR _12786_ sky130_fd_sc_hd__mux2_1
XFILLER_89_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25984_ _11287_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27723_ registers\[33\]\[11\] _10328_ _12233_ VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__mux2_1
XFILLER_24_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20058_ registers\[36\]\[48\] registers\[37\]\[48\] registers\[38\]\[48\] registers\[39\]\[48\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__mux4_1
X_24935_ _09594_ registers\[53\]\[38\] _10691_ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__mux2_1
XFILLER_86_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27654_ _12198_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__clkbuf_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24866_ _09525_ registers\[53\]\[5\] _10658_ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__mux2_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26605_ _11614_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23817_ _10077_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__clkbuf_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_224 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27585_ _12150_ VGND VGND VPWR VPWR _12162_ sky130_fd_sc_hd__buf_6
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _10627_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__clkbuf_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29324_ _09764_ registers\[22\]\[35\] _13102_ VGND VGND VPWR VPWR _13108_ sky130_fd_sc_hd__mux2_1
XFILLER_54_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26536_ _11577_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_268 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _10041_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_279 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29255_ _09662_ registers\[22\]\[2\] _13069_ VGND VGND VPWR VPWR _13072_ sky130_fd_sc_hd__mux2_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26467_ _11541_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__clkbuf_1
X_23679_ _10003_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _14540_ _14728_ _14729_ _14551_ VGND VGND VPWR VPWR _14730_ sky130_fd_sc_hd__a22o_1
X_28206_ _12488_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25418_ _10985_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__clkbuf_1
X_29186_ registers\[23\]\[43\] _13025_ _13019_ VGND VGND VPWR VPWR _13026_ sky130_fd_sc_hd__mux2_1
X_26398_ _10848_ registers\[43\]\[56\] _11498_ VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__mux2_1
XFILLER_201_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16151_ _14528_ _14661_ _14662_ _14537_ VGND VGND VPWR VPWR _14663_ sky130_fd_sc_hd__a22o_1
X_28137_ _12452_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25349_ _10949_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__clkbuf_1
X_16082_ registers\[16\]\[0\] registers\[17\]\[0\] registers\[18\]\[0\] registers\[19\]\[0\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14596_ sky130_fd_sc_hd__mux4_1
X_28068_ _11828_ registers\[31\]\[47\] _12408_ VGND VGND VPWR VPWR _12416_ sky130_fd_sc_hd__mux2_1
XFILLER_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27019_ _11862_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__clkbuf_1
X_19910_ registers\[16\]\[43\] registers\[17\]\[43\] registers\[18\]\[43\] registers\[19\]\[43\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__mux4_1
XFILLER_194_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30030_ _13423_ VGND VGND VPWR VPWR _13479_ sky130_fd_sc_hd__buf_4
X_19841_ _06525_ _06561_ _06562_ _06528_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__a22o_1
XFILLER_116_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19772_ _06495_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__buf_2
X_16984_ _15468_ _15471_ _15269_ VGND VGND VPWR VPWR _15472_ sky130_fd_sc_hd__o21ba_1
XFILLER_96_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18723_ _05469_ _05474_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31981_ clknet_leaf_21_CLK _00152_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1063 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18654_ registers\[48\]\[8\] registers\[49\]\[8\] registers\[50\]\[8\] registers\[51\]\[8\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__mux4_1
X_33720_ clknet_leaf_339_CLK _01834_ VGND VGND VPWR VPWR registers\[41\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_30932_ registers\[10\]\[29\] _12995_ _13944_ VGND VGND VPWR VPWR _13954_ sky130_fd_sc_hd__mux2_1
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_6_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17605_ registers\[12\]\[43\] registers\[13\]\[43\] registers\[14\]\[43\] registers\[15\]\[43\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__mux4_1
XFILLER_236_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30863_ _13917_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__clkbuf_1
X_18585_ registers\[52\]\[6\] registers\[53\]\[6\] registers\[54\]\[6\] registers\[55\]\[6\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__mux4_1
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33651_ clknet_leaf_348_CLK _01765_ VGND VGND VPWR VPWR registers\[42\]\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32602_ clknet_leaf_84_CLK _00716_ VGND VGND VPWR VPWR registers\[58\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17536_ registers\[4\]\[41\] registers\[5\]\[41\] registers\[6\]\[41\] registers\[7\]\[41\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__mux4_1
X_33582_ clknet_leaf_348_CLK _01696_ VGND VGND VPWR VPWR registers\[43\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30794_ _13881_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_780 _08338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32533_ clknet_leaf_74_CLK _00647_ VGND VGND VPWR VPWR registers\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_791 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35321_ clknet_leaf_310_CLK _03435_ VGND VGND VPWR VPWR registers\[16\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17467_ registers\[28\]\[39\] registers\[29\]\[39\] registers\[30\]\[39\] registers\[31\]\[39\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15942_ sky130_fd_sc_hd__mux4_1
XFILLER_60_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ _14504_ VGND VGND VPWR VPWR _14922_ sky130_fd_sc_hd__clkbuf_4
X_19206_ registers\[28\]\[23\] registers\[29\]\[23\] registers\[30\]\[23\] registers\[31\]\[23\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__mux4_1
X_32464_ clknet_leaf_176_CLK _00578_ VGND VGND VPWR VPWR registers\[60\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_35252_ clknet_leaf_417_CLK _03366_ VGND VGND VPWR VPWR registers\[17\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17398_ _15871_ _15874_ _15645_ VGND VGND VPWR VPWR _15875_ sky130_fd_sc_hd__o21ba_1
XFILLER_203_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31415_ _14208_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__clkbuf_1
X_19137_ registers\[20\]\[21\] registers\[21\]\[21\] registers\[22\]\[21\] registers\[23\]\[21\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__mux4_1
X_34203_ clknet_leaf_18_CLK _02317_ VGND VGND VPWR VPWR registers\[33\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16349_ _14527_ VGND VGND VPWR VPWR _14855_ sky130_fd_sc_hd__clkbuf_4
X_35183_ clknet_leaf_394_CLK _03297_ VGND VGND VPWR VPWR registers\[18\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_32395_ clknet_leaf_167_CLK _00509_ VGND VGND VPWR VPWR registers\[61\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34134_ clknet_leaf_122_CLK _02248_ VGND VGND VPWR VPWR registers\[34\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31346_ registers\[7\]\[33\] net27 _14168_ VGND VGND VPWR VPWR _14172_ sky130_fd_sc_hd__mux2_1
X_19068_ registers\[32\]\[20\] registers\[33\]\[20\] registers\[34\]\[20\] registers\[35\]\[20\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__mux4_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18019_ registers\[8\]\[55\] registers\[9\]\[55\] registers\[10\]\[55\] registers\[11\]\[55\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux4_2
X_34065_ clknet_leaf_134_CLK _02179_ VGND VGND VPWR VPWR registers\[35\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31277_ registers\[7\]\[0\] net1 _14135_ VGND VGND VPWR VPWR _14136_ sky130_fd_sc_hd__mux2_1
X_33016_ clknet_leaf_334_CLK _01130_ VGND VGND VPWR VPWR registers\[52\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21030_ _07338_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__clkbuf_4
X_30228_ _13583_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30159_ registers\[16\]\[47\] _13033_ _13539_ VGND VGND VPWR VPWR _13547_ sky130_fd_sc_hd__mux2_1
XFILLER_102_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34967_ clknet_leaf_99_CLK _03081_ VGND VGND VPWR VPWR registers\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_22981_ _09583_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1035 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1190 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24720_ _10586_ VGND VGND VPWR VPWR _10587_ sky130_fd_sc_hd__buf_4
X_33918_ clknet_leaf_269_CLK _02032_ VGND VGND VPWR VPWR registers\[38\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_21932_ registers\[32\]\[36\] registers\[33\]\[36\] registers\[34\]\[36\] registers\[35\]\[36\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__mux4_1
XFILLER_216_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34898_ clknet_leaf_100_CLK _03012_ VGND VGND VPWR VPWR registers\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24651_ _09582_ registers\[55\]\[32\] _10547_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__mux2_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33849_ clknet_leaf_302_CLK _01963_ VGND VGND VPWR VPWR registers\[3\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_21863_ _08505_ _08512_ _08521_ _08528_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__or4_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23602_ registers\[61\]\[18\] _09695_ _09954_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__mux2_1
XFILLER_247_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20814_ registers\[56\]\[4\] registers\[57\]\[4\] registers\[58\]\[4\] registers\[59\]\[4\]
+ _07508_ _07317_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__mux4_1
X_27370_ registers\[36\]\[37\] _10382_ _12040_ VGND VGND VPWR VPWR _12048_ sky130_fd_sc_hd__mux2_1
XFILLER_230_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24582_ _10510_ _10512_ VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__nand2_8
X_21794_ _08461_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__buf_6
XFILLER_70_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26321_ _11464_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__clkbuf_1
X_23533_ _09619_ registers\[19\]\[50\] _09925_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__mux2_1
X_35519_ clknet_leaf_297_CLK _03633_ VGND VGND VPWR VPWR registers\[13\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20745_ registers\[36\]\[2\] registers\[37\]\[2\] registers\[38\]\[2\] registers\[39\]\[2\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__mux4_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29040_ registers\[24\]\[60\] _10430_ _12860_ VGND VGND VPWR VPWR _12927_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26252_ _11428_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20676_ _07363_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__buf_4
X_23464_ _09889_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25203_ _10743_ registers\[51\]\[6\] _10865_ VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__mux2_1
X_22415_ _08958_ _09063_ _09064_ _08961_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__a22o_1
XFILLER_137_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26183_ _10768_ registers\[44\]\[18\] _11383_ VGND VGND VPWR VPWR _11392_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23395_ registers\[39\]\[50\] _09797_ _09851_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__mux2_1
XFILLER_164_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25134_ net41 VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__buf_2
X_22346_ registers\[16\]\[47\] registers\[17\]\[47\] registers\[18\]\[47\] registers\[19\]\[47\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__mux4_1
XFILLER_100_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22277_ _08761_ _08929_ _08930_ _08764_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__a22o_1
X_29942_ registers\[17\]\[8\] _12951_ _13424_ VGND VGND VPWR VPWR _13433_ sky130_fd_sc_hd__mux2_1
X_25065_ _10780_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
X_24016_ _10160_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__buf_4
X_21228_ registers\[44\]\[16\] registers\[45\]\[16\] registers\[46\]\[16\] registers\[47\]\[16\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29873_ _13396_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28824_ _11774_ registers\[25\]\[21\] _12812_ VGND VGND VPWR VPWR _12814_ sky130_fd_sc_hd__mux2_1
X_21159_ registers\[40\]\[14\] registers\[41\]\[14\] registers\[42\]\[14\] registers\[43\]\[14\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__mux4_1
X_28755_ _12777_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25967_ _11278_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27706_ registers\[33\]\[3\] _10311_ _12222_ VGND VGND VPWR VPWR _12226_ sky130_fd_sc_hd__mux2_1
XFILLER_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24918_ _10657_ VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__clkbuf_8
X_28686_ _12718_ VGND VGND VPWR VPWR _12741_ sky130_fd_sc_hd__buf_4
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25898_ _11242_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27637_ _12189_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__clkbuf_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24849_ _10654_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18370_ net81 net82 VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__or2_4
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27568_ _12153_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__clkbuf_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17321_ _15796_ _15799_ _15631_ VGND VGND VPWR VPWR _15800_ sky130_fd_sc_hd__o21ba_1
X_29307_ _09747_ registers\[22\]\[27\] _13091_ VGND VGND VPWR VPWR _13099_ sky130_fd_sc_hd__mux2_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26519_ _11568_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27499_ _11801_ registers\[35\]\[34\] _12111_ VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__mux2_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29238_ registers\[23\]\[60\] _13060_ _12934_ VGND VGND VPWR VPWR _13061_ sky130_fd_sc_hd__mux2_1
X_17252_ registers\[12\]\[33\] registers\[13\]\[33\] registers\[14\]\[33\] registers\[15\]\[33\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15733_ sky130_fd_sc_hd__mux4_1
XFILLER_35_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16203_ _14710_ _14713_ _14614_ VGND VGND VPWR VPWR _14714_ sky130_fd_sc_hd__o21ba_1
XFILLER_168_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17183_ registers\[4\]\[31\] registers\[5\]\[31\] registers\[6\]\[31\] registers\[7\]\[31\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15666_ sky130_fd_sc_hd__mux4_1
XFILLER_31_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29169_ net32 VGND VGND VPWR VPWR _13014_ sky130_fd_sc_hd__buf_2
X_31200_ registers\[8\]\[28\] net21 _14086_ VGND VGND VPWR VPWR _14095_ sky130_fd_sc_hd__mux2_1
X_16134_ _14625_ _14632_ _14639_ _14646_ VGND VGND VPWR VPWR _14647_ sky130_fd_sc_hd__or4_2
X_32180_ clknet_leaf_484_CLK _00294_ VGND VGND VPWR VPWR registers\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_31131_ _14058_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__clkbuf_1
X_16065_ _14578_ VGND VGND VPWR VPWR _14579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31062_ _14022_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30013_ _13470_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19824_ _06542_ _06545_ _06504_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__o21ba_1
XFILLER_190_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35870_ clknet_leaf_480_CLK _03984_ VGND VGND VPWR VPWR registers\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34821_ clknet_leaf_225_CLK _02935_ VGND VGND VPWR VPWR registers\[24\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19755_ _06441_ _06477_ _06478_ _06445_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__a22o_1
X_16967_ _15144_ _15454_ _15455_ _15147_ VGND VGND VPWR VPWR _15456_ sky130_fd_sc_hd__a22o_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18706_ registers\[16\]\[9\] registers\[17\]\[9\] registers\[18\]\[9\] registers\[19\]\[9\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__mux4_1
X_34752_ clknet_leaf_226_CLK _02866_ VGND VGND VPWR VPWR registers\[25\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16898_ _14520_ VGND VGND VPWR VPWR _15389_ sky130_fd_sc_hd__buf_4
X_31964_ clknet_leaf_4_CLK _00133_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
X_19686_ registers\[0\]\[37\] registers\[1\]\[37\] registers\[2\]\[37\] registers\[3\]\[37\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__mux4_1
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33703_ clknet_leaf_430_CLK _01817_ VGND VGND VPWR VPWR registers\[41\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_18637_ registers\[20\]\[7\] registers\[21\]\[7\] registers\[22\]\[7\] registers\[23\]\[7\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__mux4_1
X_30915_ _13945_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__clkbuf_1
X_34683_ clknet_leaf_183_CLK _02797_ VGND VGND VPWR VPWR registers\[26\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31895_ _14460_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30846_ _09802_ registers\[11\]\[52\] _13906_ VGND VGND VPWR VPWR _13909_ sky130_fd_sc_hd__mux2_1
XFILLER_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33634_ clknet_leaf_55_CLK _01748_ VGND VGND VPWR VPWR registers\[42\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18568_ _05150_ _05324_ _05325_ _05160_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__a22o_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17519_ registers\[32\]\[41\] registers\[33\]\[41\] registers\[34\]\[41\] registers\[35\]\[41\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__mux4_1
X_18499_ _05137_ _05257_ _05258_ _05147_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__a22o_1
X_30777_ _13872_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__clkbuf_1
X_33565_ clknet_leaf_28_CLK _01679_ VGND VGND VPWR VPWR registers\[43\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20530_ registers\[0\]\[62\] registers\[1\]\[62\] registers\[2\]\[62\] registers\[3\]\[62\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__mux4_1
X_35304_ clknet_leaf_404_CLK _03418_ VGND VGND VPWR VPWR registers\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_32516_ clknet_leaf_201_CLK _00630_ VGND VGND VPWR VPWR registers\[60\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_33496_ clknet_leaf_34_CLK _01610_ VGND VGND VPWR VPWR registers\[44\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20461_ _07160_ _07163_ _05073_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__o21ba_1
X_32447_ clknet_leaf_306_CLK _00561_ VGND VGND VPWR VPWR registers\[29\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_35235_ clknet_leaf_474_CLK _03349_ VGND VGND VPWR VPWR registers\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22200_ registers\[8\]\[43\] registers\[9\]\[43\] registers\[10\]\[43\] registers\[11\]\[43\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__mux4_1
X_23180_ registers\[9\]\[8\] _09674_ _09709_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__mux2_1
X_20392_ _07094_ _07097_ _06880_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__o21ba_1
X_32378_ clknet_leaf_287_CLK _00492_ VGND VGND VPWR VPWR registers\[61\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35166_ clknet_leaf_1_CLK _03280_ VGND VGND VPWR VPWR registers\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22131_ _08785_ _08788_ _08748_ _08749_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__o211a_1
X_34117_ clknet_leaf_246_CLK _02231_ VGND VGND VPWR VPWR registers\[35\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_31329_ registers\[7\]\[25\] net18 _14157_ VGND VGND VPWR VPWR _14163_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35097_ clknet_leaf_11_CLK _03211_ VGND VGND VPWR VPWR registers\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xoutput220 net220 VGND VGND VPWR VPWR D3[11] sky130_fd_sc_hd__buf_2
Xoutput231 net231 VGND VGND VPWR VPWR D3[21] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR D3[31] sky130_fd_sc_hd__buf_2
XTAP_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput253 net253 VGND VGND VPWR VPWR D3[41] sky130_fd_sc_hd__buf_2
X_22062_ _08615_ _08720_ _08721_ _08618_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__a22o_1
XTAP_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34048_ clknet_leaf_258_CLK _02162_ VGND VGND VPWR VPWR registers\[36\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput264 net264 VGND VGND VPWR VPWR D3[51] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR D3[61] sky130_fd_sc_hd__buf_2
Xclkbuf_6_3__f_CLK clknet_5_1_0_CLK VGND VGND VPWR VPWR clknet_6_3__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21013_ _07702_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
XTAP_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26870_ _11761_ registers\[3\]\[15\] _11751_ VGND VGND VPWR VPWR _11762_ sky130_fd_sc_hd__mux2_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25821_ _11201_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35999_ clknet_leaf_46_CLK _04113_ VGND VGND VPWR VPWR registers\[63\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28540_ _12664_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__clkbuf_1
X_25752_ _11165_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22964_ _09571_ registers\[62\]\[27\] _09557_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24703_ _09634_ registers\[55\]\[57\] _10569_ VGND VGND VPWR VPWR _10577_ sky130_fd_sc_hd__mux2_1
XFILLER_243_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28471_ _11826_ registers\[28\]\[46\] _12621_ VGND VGND VPWR VPWR _12628_ sky130_fd_sc_hd__mux2_1
X_21915_ registers\[8\]\[35\] registers\[9\]\[35\] registers\[10\]\[35\] registers\[11\]\[35\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__mux4_1
X_25683_ registers\[48\]\[38\] _10384_ _11119_ VGND VGND VPWR VPWR _11128_ sky130_fd_sc_hd__mux2_1
X_22895_ net56 VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27422_ registers\[36\]\[62\] _10434_ _12006_ VGND VGND VPWR VPWR _12075_ sky130_fd_sc_hd__mux2_1
XFILLER_243_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24634_ _09565_ registers\[55\]\[24\] _10536_ VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__mux2_1
XFILLER_130_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21846_ _08508_ _08511_ _08405_ _08406_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__o211a_1
XFILLER_224_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27353_ registers\[36\]\[29\] _10365_ _12029_ VGND VGND VPWR VPWR _12039_ sky130_fd_sc_hd__mux2_1
XFILLER_230_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24565_ _09634_ registers\[56\]\[57\] _10495_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__mux2_1
XFILLER_24_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21777_ _08334_ _08443_ _08444_ _08338_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__a22o_1
XFILLER_19_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26304_ _10754_ registers\[43\]\[11\] _11454_ VGND VGND VPWR VPWR _11456_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23516_ _09603_ registers\[19\]\[42\] _09914_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__mux2_1
X_27284_ _12002_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__clkbuf_1
X_20728_ registers\[16\]\[1\] registers\[17\]\[1\] registers\[18\]\[1\] registers\[19\]\[1\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__mux4_1
XFILLER_157_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24496_ _09565_ registers\[56\]\[24\] _10462_ VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__mux2_1
XFILLER_211_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29023_ _12918_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26235_ _11419_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23447_ _09880_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__clkbuf_1
X_20659_ _07280_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__buf_12
XFILLER_17_1092 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26166_ _11371_ VGND VGND VPWR VPWR _11383_ sky130_fd_sc_hd__buf_4
X_23378_ registers\[39\]\[42\] _09780_ _09840_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__mux2_1
XFILLER_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25117_ _10814_ registers\[52\]\[40\] _10815_ VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__mux2_1
X_22329_ _08812_ _08977_ _08980_ _08815_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__a22o_1
XFILLER_87_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26097_ _10817_ registers\[45\]\[41\] _11345_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29925_ _13423_ VGND VGND VPWR VPWR _13424_ sky130_fd_sc_hd__buf_6
X_25048_ _10768_ registers\[52\]\[18\] _10752_ VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__mux2_1
XFILLER_140_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17870_ _04646_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_2
XFILLER_151_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29856_ registers\[18\]\[31\] _13000_ _13386_ VGND VGND VPWR VPWR _13388_ sky130_fd_sc_hd__mux2_1
XFILLER_66_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28807_ _11757_ registers\[25\]\[13\] _12801_ VGND VGND VPWR VPWR _12805_ sky130_fd_sc_hd__mux2_1
X_16821_ _15198_ _15312_ _15313_ _15204_ VGND VGND VPWR VPWR _15314_ sky130_fd_sc_hd__a22o_1
XFILLER_232_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29787_ registers\[1\]\[63\] _13066_ _13281_ VGND VGND VPWR VPWR _13351_ sky130_fd_sc_hd__mux2_1
X_26999_ net53 VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__buf_4
XFILLER_19_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19540_ registers\[56\]\[33\] registers\[57\]\[33\] registers\[58\]\[33\] registers\[59\]\[33\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__mux4_1
X_16752_ registers\[0\]\[19\] registers\[1\]\[19\] registers\[2\]\[19\] registers\[3\]\[19\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15247_ sky130_fd_sc_hd__mux4_1
XFILLER_4_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28738_ _12768_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16683_ registers\[4\]\[17\] registers\[5\]\[17\] registers\[6\]\[17\] registers\[7\]\[17\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15180_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28669_ _12732_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__clkbuf_1
X_19471_ _06199_ _06202_ _06161_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__o21ba_1
XFILLER_234_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30700_ registers\[12\]\[47\] _13033_ _13824_ VGND VGND VPWR VPWR _13832_ sky130_fd_sc_hd__mux2_1
XFILLER_222_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18422_ _05107_ _05182_ _05183_ _05117_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__a22o_1
X_31680_ _09867_ _09940_ VGND VGND VPWR VPWR _14347_ sky130_fd_sc_hd__nor2_8
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18353_ _05048_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__buf_12
X_30631_ registers\[12\]\[14\] _12964_ _13791_ VGND VGND VPWR VPWR _13796_ sky130_fd_sc_hd__mux2_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_230_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_230_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _15684_ _15781_ _15782_ _15687_ VGND VGND VPWR VPWR _15783_ sky130_fd_sc_hd__a22o_1
X_33350_ clknet_leaf_254_CLK _01464_ VGND VGND VPWR VPWR registers\[47\]\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ registers\[40\]\[0\] registers\[41\]\[0\] registers\[42\]\[0\] registers\[43\]\[0\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__mux4_1
X_30562_ _13759_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32301_ clknet_leaf_397_CLK _00415_ VGND VGND VPWR VPWR registers\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17235_ _15677_ _15714_ _15715_ _15682_ VGND VGND VPWR VPWR _15716_ sky130_fd_sc_hd__a22o_1
X_33281_ clknet_leaf_270_CLK _01395_ VGND VGND VPWR VPWR registers\[48\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30493_ _13723_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32232_ clknet_leaf_144_CLK _00346_ VGND VGND VPWR VPWR registers\[9\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_35020_ clknet_leaf_143_CLK _03134_ VGND VGND VPWR VPWR registers\[21\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17166_ registers\[32\]\[31\] registers\[33\]\[31\] registers\[34\]\[31\] registers\[35\]\[31\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15649_ sky130_fd_sc_hd__mux4_1
XFILLER_122_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16117_ registers\[52\]\[1\] registers\[53\]\[1\] registers\[54\]\[1\] registers\[55\]\[1\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14630_ sky130_fd_sc_hd__mux4_1
XFILLER_116_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32163_ clknet_leaf_440_CLK _00277_ VGND VGND VPWR VPWR registers\[39\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17097_ registers\[56\]\[29\] registers\[57\]\[29\] registers\[58\]\[29\] registers\[59\]\[29\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15582_ sky130_fd_sc_hd__mux4_1
XFILLER_196_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31114_ registers\[0\]\[51\] _13042_ _14048_ VGND VGND VPWR VPWR _14050_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16048_ _14529_ VGND VGND VPWR VPWR _14562_ sky130_fd_sc_hd__buf_12
X_32094_ clknet_leaf_485_CLK _00007_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_297_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_297_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35922_ clknet_leaf_77_CLK _04036_ VGND VGND VPWR VPWR registers\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_31045_ _14013_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19807_ _05059_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__clkbuf_4
X_35853_ clknet_leaf_144_CLK _03967_ VGND VGND VPWR VPWR registers\[8\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_17999_ registers\[28\]\[54\] registers\[29\]\[54\] registers\[30\]\[54\] registers\[31\]\[54\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__mux4_1
X_34804_ clknet_leaf_414_CLK _02918_ VGND VGND VPWR VPWR registers\[24\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_19738_ _06459_ _06462_ _06194_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__o21ba_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35784_ clknet_leaf_217_CLK _03898_ VGND VGND VPWR VPWR registers\[0\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32996_ clknet_leaf_442_CLK _01110_ VGND VGND VPWR VPWR registers\[52\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_231_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34735_ clknet_leaf_386_CLK _02849_ VGND VGND VPWR VPWR registers\[25\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_31947_ _14487_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__clkbuf_1
X_19669_ registers\[40\]\[37\] registers\[41\]\[37\] registers\[42\]\[37\] registers\[43\]\[37\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__mux4_1
XFILLER_20_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21700_ registers\[60\]\[29\] registers\[61\]\[29\] registers\[62\]\[29\] registers\[63\]\[29\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__mux4_1
XFILLER_240_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22680_ registers\[0\]\[57\] registers\[1\]\[57\] registers\[2\]\[57\] registers\[3\]\[57\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__mux4_1
XFILLER_240_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34666_ clknet_leaf_452_CLK _02780_ VGND VGND VPWR VPWR registers\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_31878_ _14451_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33617_ clknet_leaf_129_CLK _01731_ VGND VGND VPWR VPWR registers\[42\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_21631_ _08299_ _08302_ _08062_ _08063_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__o211a_1
XFILLER_209_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30829_ _09784_ registers\[11\]\[44\] _13895_ VGND VGND VPWR VPWR _13900_ sky130_fd_sc_hd__mux2_1
X_34597_ clknet_leaf_445_CLK _02711_ VGND VGND VPWR VPWR registers\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_221_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_221_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_205_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24350_ _10375_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
X_33548_ clknet_leaf_176_CLK _01662_ VGND VGND VPWR VPWR registers\[44\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_21562_ registers\[8\]\[25\] registers\[9\]\[25\] registers\[10\]\[25\] registers\[11\]\[25\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__mux4_1
XFILLER_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23301_ registers\[9\]\[49\] _09795_ _09776_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__mux2_1
XFILLER_138_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20513_ _07193_ _07200_ _07207_ _07214_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__or4_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24281_ registers\[57\]\[11\] _10328_ _10326_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__mux2_1
X_21493_ _08165_ _08168_ _08062_ _08063_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__o211a_1
X_33479_ clknet_leaf_250_CLK _01593_ VGND VGND VPWR VPWR registers\[45\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26020_ _11306_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20444_ _05060_ _07146_ _07147_ _05066_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__a22o_1
X_35218_ clknet_leaf_101_CLK _03332_ VGND VGND VPWR VPWR registers\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_23232_ registers\[9\]\[28\] _09749_ _09735_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__mux2_1
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36198_ clknet_leaf_98_CLK _00080_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35149_ clknet_leaf_147_CLK _03263_ VGND VGND VPWR VPWR registers\[1\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_23163_ registers\[9\]\[1\] _09660_ _09709_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__mux2_1
X_20375_ registers\[60\]\[57\] registers\[61\]\[57\] registers\[62\]\[57\] registers\[63\]\[57\]
+ _06991_ _06785_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__mux4_1
XTAP_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22114_ _07398_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__clkbuf_4
XTAP_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23094_ registers\[39\]\[2\] _09662_ _09658_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__mux2_1
X_27971_ _12365_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__clkbuf_1
XTAP_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_288_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_288_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26922_ net26 VGND VGND VPWR VPWR _11797_ sky130_fd_sc_hd__clkbuf_4
X_29710_ registers\[1\]\[26\] _12989_ _13304_ VGND VGND VPWR VPWR _13311_ sky130_fd_sc_hd__mux2_1
X_22045_ _08462_ _08701_ _08704_ _08467_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__a22o_1
XTAP_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29641_ _13274_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__clkbuf_1
XTAP_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26853_ net2 VGND VGND VPWR VPWR _11750_ sky130_fd_sc_hd__clkbuf_4
XFILLER_216_1399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25804_ _10793_ registers\[47\]\[30\] _11192_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__mux2_1
XFILLER_217_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29572_ _13238_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__clkbuf_1
X_26784_ registers\[40\]\[46\] _10401_ _11702_ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23996_ _09535_ registers\[5\]\[10\] _10172_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__mux2_1
XFILLER_229_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28523_ _12655_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25735_ registers\[48\]\[63\] _10436_ _11085_ VGND VGND VPWR VPWR _11155_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22947_ _09560_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_460_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_460_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28454_ _11809_ registers\[28\]\[38\] _12610_ VGND VGND VPWR VPWR _12619_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25666_ _11085_ VGND VGND VPWR VPWR _11119_ sky130_fd_sc_hd__buf_4
X_22878_ _09511_ net83 _09512_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__or3b_1
XFILLER_231_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27405_ _12066_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__clkbuf_1
X_24617_ _09548_ registers\[55\]\[16\] _10525_ VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__mux2_1
X_28385_ _11740_ registers\[28\]\[5\] _12577_ VGND VGND VPWR VPWR _12583_ sky130_fd_sc_hd__mux2_1
X_21829_ _08423_ _08494_ _08495_ _08428_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__a22o_1
X_25597_ registers\[4\]\[63\] _10436_ _11011_ VGND VGND VPWR VPWR _11081_ sky130_fd_sc_hd__mux2_1
XFILLER_169_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_212_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_212_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27336_ _12030_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_1
X_24548_ _09617_ registers\[56\]\[49\] _10484_ VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27267_ _11839_ registers\[37\]\[52\] _11991_ VGND VGND VPWR VPWR _11994_ sky130_fd_sc_hd__mux2_1
XFILLER_8_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24479_ _09548_ registers\[56\]\[16\] _10451_ VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__mux2_1
X_29006_ _12909_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__clkbuf_1
X_17020_ _14571_ VGND VGND VPWR VPWR _15507_ sky130_fd_sc_hd__buf_6
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26218_ _11410_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27198_ _11957_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_15_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_15_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26149_ _11374_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18971_ _05711_ _05716_ _05475_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__o21ba_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_279_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_279_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1701 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29908_ registers\[18\]\[56\] _13052_ _13408_ VGND VGND VPWR VPWR _13415_ sky130_fd_sc_hd__mux2_1
X_17922_ registers\[0\]\[52\] registers\[1\]\[52\] registers\[2\]\[52\] registers\[3\]\[52\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux4_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1712 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1723 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1734 _00180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1745 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1756 _07315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17853_ _14584_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__buf_2
XANTENNA_1767 _08943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29839_ registers\[18\]\[23\] _12983_ _13375_ VGND VGND VPWR VPWR _13379_ sky130_fd_sc_hd__mux2_1
XFILLER_66_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1778 _12006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1789 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16804_ _14607_ VGND VGND VPWR VPWR _15298_ sky130_fd_sc_hd__clkbuf_4
X_32850_ clknet_leaf_64_CLK _00964_ VGND VGND VPWR VPWR registers\[54\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17784_ _04557_ _04562_ _15974_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__o21ba_1
XFILLER_82_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31801_ registers\[59\]\[57\] net53 _14403_ VGND VGND VPWR VPWR _14411_ sky130_fd_sc_hd__mux2_1
X_19523_ registers\[16\]\[32\] registers\[17\]\[32\] registers\[18\]\[32\] registers\[19\]\[32\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__mux4_1
XFILLER_47_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16735_ registers\[40\]\[19\] registers\[41\]\[19\] registers\[42\]\[19\] registers\[43\]\[19\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15230_ sky130_fd_sc_hd__mux4_1
X_32781_ clknet_leaf_140_CLK _00895_ VGND VGND VPWR VPWR registers\[56\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_451_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_451_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34520_ clknet_leaf_15_CLK _02634_ VGND VGND VPWR VPWR registers\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_19454_ _05149_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__clkbuf_4
X_31732_ registers\[59\]\[24\] net17 _14370_ VGND VGND VPWR VPWR _14375_ sky130_fd_sc_hd__mux2_1
X_16666_ registers\[44\]\[17\] registers\[45\]\[17\] registers\[46\]\[17\] registers\[47\]\[17\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15163_ sky130_fd_sc_hd__mux4_1
XFILLER_234_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18405_ registers\[32\]\[1\] registers\[33\]\[1\] registers\[34\]\[1\] registers\[35\]\[1\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__mux4_1
X_34451_ clknet_leaf_105_CLK _02565_ VGND VGND VPWR VPWR registers\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31663_ _14338_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__clkbuf_1
X_19385_ _06116_ _06119_ _05851_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__o21ba_1
XFILLER_50_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16597_ registers\[36\]\[15\] registers\[37\]\[15\] registers\[38\]\[15\] registers\[39\]\[15\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _15096_ sky130_fd_sc_hd__mux4_1
XFILLER_61_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_203_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_203_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33402_ clknet_leaf_279_CLK _01516_ VGND VGND VPWR VPWR registers\[46\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18336_ registers\[52\]\[0\] registers\[53\]\[0\] registers\[54\]\[0\] registers\[55\]\[0\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__mux4_1
X_30614_ registers\[12\]\[6\] _12947_ _13780_ VGND VGND VPWR VPWR _13787_ sky130_fd_sc_hd__mux2_1
XFILLER_148_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34382_ clknet_leaf_109_CLK _02496_ VGND VGND VPWR VPWR registers\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31594_ _14302_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36121_ clknet_leaf_35_CLK _04235_ VGND VGND VPWR VPWR registers\[49\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18267_ registers\[16\]\[63\] registers\[17\]\[63\] registers\[18\]\[63\] registers\[19\]\[63\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__mux4_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30545_ _13750_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__clkbuf_1
X_33333_ clknet_leaf_344_CLK _01447_ VGND VGND VPWR VPWR registers\[47\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36052_ clknet_leaf_71_CLK _04166_ VGND VGND VPWR VPWR registers\[59\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17218_ registers\[12\]\[32\] registers\[13\]\[32\] registers\[14\]\[32\] registers\[15\]\[32\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15700_ sky130_fd_sc_hd__mux4_1
X_18198_ _04960_ _04963_ _14553_ _14555_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__o211a_1
X_30476_ _13714_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33264_ clknet_leaf_366_CLK _01378_ VGND VGND VPWR VPWR registers\[48\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_35003_ clknet_leaf_307_CLK _03117_ VGND VGND VPWR VPWR registers\[21\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_17149_ _14587_ VGND VGND VPWR VPWR _15633_ sky130_fd_sc_hd__clkbuf_4
X_32215_ clknet_leaf_435_CLK _00329_ VGND VGND VPWR VPWR registers\[39\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_33195_ clknet_leaf_402_CLK _01309_ VGND VGND VPWR VPWR registers\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_16__f_CLK clknet_5_8_0_CLK VGND VGND VPWR VPWR clknet_6_16__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_32146_ clknet_leaf_119_CLK _00260_ VGND VGND VPWR VPWR registers\[39\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20160_ _05059_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_131_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32077_ clknet_leaf_167_CLK _00255_ VGND VGND VPWR VPWR registers\[62\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20091_ _06802_ _06805_ _06537_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__o21ba_1
XFILLER_170_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35905_ clknet_leaf_234_CLK _04019_ VGND VGND VPWR VPWR registers\[7\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_31028_ registers\[0\]\[10\] _12955_ _14004_ VGND VGND VPWR VPWR _14005_ sky130_fd_sc_hd__mux2_1
XFILLER_44_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23850_ _10095_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
X_35836_ clknet_leaf_300_CLK _03950_ VGND VGND VPWR VPWR registers\[8\]\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22801_ _07276_ _09437_ _09438_ _07286_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__a22o_1
XFILLER_66_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35767_ clknet_leaf_314_CLK _03881_ VGND VGND VPWR VPWR registers\[0\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_23781_ _10058_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_609 _05111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32979_ clknet_leaf_72_CLK _01093_ VGND VGND VPWR VPWR registers\[52\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_20993_ _07640_ _07681_ _07682_ _07646_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a22o_1
XFILLER_66_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25520_ registers\[4\]\[26\] _10359_ _11034_ VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_442_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_442_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_246_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22732_ registers\[56\]\[59\] registers\[57\]\[59\] registers\[58\]\[59\] registers\[59\]\[59\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34718_ clknet_leaf_3_CLK _02832_ VGND VGND VPWR VPWR registers\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35698_ clknet_leaf_382_CLK _03812_ VGND VGND VPWR VPWR registers\[10\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_25451_ _11002_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22663_ _09284_ _09291_ _09298_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__or4_4
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34649_ clknet_leaf_21_CLK _02763_ VGND VGND VPWR VPWR registers\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24402_ registers\[57\]\[50\] _10409_ _10410_ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28170_ _11795_ registers\[30\]\[31\] _12468_ VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__mux2_1
X_21614_ _08257_ _08266_ _08277_ _08286_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__or4_4
X_25382_ _10966_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_1
X_22594_ _07347_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__buf_6
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27121_ _11828_ registers\[38\]\[47\] _11909_ VGND VGND VPWR VPWR _11917_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24333_ registers\[57\]\[28\] _10363_ _10347_ VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__mux2_1
XFILLER_107_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21545_ _08219_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27052_ _11759_ registers\[38\]\[14\] _11876_ VGND VGND VPWR VPWR _11881_ sky130_fd_sc_hd__mux2_1
X_24264_ net61 VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__buf_4
XFILLER_181_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21476_ _08080_ _08151_ _08152_ _08085_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__a22o_1
XFILLER_193_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26003_ _10858_ registers\[46\]\[61\] _11229_ VGND VGND VPWR VPWR _11297_ sky130_fd_sc_hd__mux2_1
X_23215_ registers\[9\]\[23\] _09730_ _09735_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__mux2_1
X_20427_ _06912_ _07129_ _07130_ _06917_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24195_ _09598_ registers\[58\]\[40\] _10277_ VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__mux2_1
XFILLER_135_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23146_ registers\[39\]\[19\] _09697_ _09679_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__mux2_1
X_20358_ _06868_ _07063_ _07064_ _06871_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__a22o_1
XTAP_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1008 _11853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27954_ registers\[32\]\[57\] _10424_ _12348_ VGND VGND VPWR VPWR _12356_ sky130_fd_sc_hd__mux2_1
X_20289_ _06717_ _06996_ _06997_ _06720_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__a22o_1
XANTENNA_1019 _12434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23077_ net1 VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__buf_4
XFILLER_62_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26905_ _11785_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_1
X_22028_ _07363_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__buf_4
XTAP_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27885_ registers\[32\]\[24\] _10355_ _12315_ VGND VGND VPWR VPWR _12320_ sky130_fd_sc_hd__mux2_1
XFILLER_212_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29624_ _13265_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26836_ _11738_ registers\[3\]\[4\] _11730_ VGND VGND VPWR VPWR _11739_ sky130_fd_sc_hd__mux2_1
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29555_ _13229_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26767_ registers\[40\]\[38\] _10384_ _11691_ VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__mux2_1
X_23979_ _09519_ registers\[5\]\[2\] _10161_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__mux2_1
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16520_ _14603_ VGND VGND VPWR VPWR _15022_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_433_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_433_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28506_ _11861_ registers\[28\]\[63\] _12576_ VGND VGND VPWR VPWR _12646_ sky130_fd_sc_hd__mux2_1
X_25718_ _11146_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26698_ registers\[40\]\[5\] _10315_ _11658_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__mux2_1
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29486_ _09793_ registers\[21\]\[48\] _13184_ VGND VGND VPWR VPWR _13193_ sky130_fd_sc_hd__mux2_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16451_ _14607_ VGND VGND VPWR VPWR _14955_ sky130_fd_sc_hd__buf_4
XFILLER_232_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28437_ _12576_ VGND VGND VPWR VPWR _12610_ sky130_fd_sc_hd__buf_4
X_25649_ _11110_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19170_ registers\[16\]\[22\] registers\[17\]\[22\] registers\[18\]\[22\] registers\[19\]\[22\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__mux4_1
X_28368_ _12573_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__clkbuf_1
X_16382_ registers\[40\]\[9\] registers\[41\]\[9\] registers\[42\]\[9\] registers\[43\]\[9\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14887_ sky130_fd_sc_hd__mux4_1
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18121_ _04637_ _04888_ _04889_ _04642_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a22o_1
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27319_ _12021_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__clkbuf_1
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28299_ _12537_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30330_ _13636_ _10585_ VGND VGND VPWR VPWR _13637_ sky130_fd_sc_hd__nand2_8
X_18052_ registers\[12\]\[56\] registers\[13\]\[56\] registers\[14\]\[56\] registers\[15\]\[56\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__mux4_1
XFILLER_240_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17003_ _15487_ _15488_ _15489_ _15490_ VGND VGND VPWR VPWR _15491_ sky130_fd_sc_hd__a22o_1
XFILLER_201_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30261_ registers\[15\]\[31\] _13000_ _13599_ VGND VGND VPWR VPWR _13601_ sky130_fd_sc_hd__mux2_1
XANTENNA_5 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32000_ clknet_leaf_27_CLK _00173_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30192_ registers\[16\]\[63\] _13066_ _13494_ VGND VGND VPWR VPWR _13564_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18954_ _05143_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__buf_4
XFILLER_79_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1520 _08841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1531 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17905_ registers\[32\]\[52\] registers\[33\]\[52\] registers\[34\]\[52\] registers\[35\]\[52\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__mux4_1
XANTENNA_1542 _10232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1553 _11513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33951_ clknet_leaf_16_CLK _02065_ VGND VGND VPWR VPWR registers\[37\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18885_ registers\[16\]\[14\] registers\[17\]\[14\] registers\[18\]\[14\] registers\[19\]\[14\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__mux4_1
XTAP_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1564 _11845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1575 _13637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1586 _14493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32902_ clknet_leaf_194_CLK _01016_ VGND VGND VPWR VPWR registers\[54\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_17836_ registers\[56\]\[50\] registers\[57\]\[50\] registers\[58\]\[50\] registers\[59\]\[50\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__mux4_1
XANTENNA_1597 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33882_ clknet_leaf_22_CLK _01996_ VGND VGND VPWR VPWR registers\[38\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_35621_ clknet_leaf_465_CLK _03735_ VGND VGND VPWR VPWR registers\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_32833_ clknet_leaf_201_CLK _00947_ VGND VGND VPWR VPWR registers\[55\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17767_ _14499_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_424_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_424_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_208_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19506_ _06233_ _06234_ _06235_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__a22o_1
X_16718_ registers\[0\]\[18\] registers\[1\]\[18\] registers\[2\]\[18\] registers\[3\]\[18\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15214_ sky130_fd_sc_hd__mux4_1
X_35552_ clknet_leaf_483_CLK _03666_ VGND VGND VPWR VPWR registers\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32764_ clknet_leaf_289_CLK _00878_ VGND VGND VPWR VPWR registers\[56\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_17698_ _15892_ _04475_ _04478_ _15896_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a22o_1
XFILLER_207_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34503_ clknet_leaf_216_CLK _02617_ VGND VGND VPWR VPWR registers\[2\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_19437_ _05104_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__clkbuf_4
X_31715_ registers\[59\]\[16\] net8 _14359_ VGND VGND VPWR VPWR _14366_ sky130_fd_sc_hd__mux2_1
X_16649_ _14581_ VGND VGND VPWR VPWR _15147_ sky130_fd_sc_hd__clkbuf_4
X_35483_ clknet_leaf_477_CLK _03597_ VGND VGND VPWR VPWR registers\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32695_ clknet_leaf_334_CLK _00809_ VGND VGND VPWR VPWR registers\[57\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34434_ clknet_leaf_221_CLK _02548_ VGND VGND VPWR VPWR registers\[30\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31646_ _14329_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__clkbuf_1
X_19368_ _06098_ _06100_ _06101_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a22o_1
XFILLER_241_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18319_ registers\[56\]\[0\] registers\[57\]\[0\] registers\[58\]\[0\] registers\[59\]\[0\]
+ _05079_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__mux4_1
XFILLER_176_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34365_ clknet_leaf_182_CLK _02479_ VGND VGND VPWR VPWR registers\[31\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31577_ _14293_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__clkbuf_1
X_19299_ _05059_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_241_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36104_ clknet_leaf_193_CLK _04218_ VGND VGND VPWR VPWR registers\[59\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33316_ clknet_leaf_62_CLK _01430_ VGND VGND VPWR VPWR registers\[47\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21330_ registers\[20\]\[18\] registers\[21\]\[18\] registers\[22\]\[18\] registers\[23\]\[18\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__mux4_1
XFILLER_135_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30528_ _13741_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34296_ clknet_leaf_338_CLK _02410_ VGND VGND VPWR VPWR registers\[32\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36035_ clknet_leaf_293_CLK _04149_ VGND VGND VPWR VPWR registers\[63\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30459_ _09821_ registers\[14\]\[61\] _13637_ VGND VGND VPWR VPWR _13705_ sky130_fd_sc_hd__mux2_1
X_33247_ clknet_leaf_35_CLK _01361_ VGND VGND VPWR VPWR registers\[48\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_21261_ _07914_ _07923_ _07934_ _07943_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__or4_1
XFILLER_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23000_ net33 VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__buf_2
X_20212_ _06919_ _06920_ _06921_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__a22o_1
XFILLER_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21192_ _07876_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33178_ clknet_leaf_13_CLK _01292_ VGND VGND VPWR VPWR registers\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20143_ _05104_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32129_ clknet_leaf_397_CLK _00046_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20074_ _06784_ _06786_ _06787_ _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__a22o_1
XFILLER_135_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24951_ _10708_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__clkbuf_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23902_ _09577_ registers\[60\]\[30\] _10122_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__mux2_1
X_27670_ registers\[34\]\[50\] _10409_ _12206_ VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__mux2_1
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24882_ _10672_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1096 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26621_ _10800_ registers\[41\]\[33\] _11619_ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23833_ _10085_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__clkbuf_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35819_ clknet_leaf_398_CLK _03933_ VGND VGND VPWR VPWR registers\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_406 _00098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_417 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_415_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_415_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26552_ _10728_ registers\[41\]\[0\] _11586_ VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__mux2_1
X_29340_ _13116_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__clkbuf_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_428 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23764_ _10049_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ registers\[28\]\[8\] registers\[29\]\[8\] registers\[30\]\[8\] registers\[31\]\[8\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__mux4_1
XANTENNA_439 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25503_ registers\[4\]\[18\] _10342_ _11023_ VGND VGND VPWR VPWR _11032_ sky130_fd_sc_hd__mux2_1
X_22715_ _09352_ _09355_ _09102_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__o21ba_1
XFILLER_199_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29271_ _13068_ VGND VGND VPWR VPWR _13080_ sky130_fd_sc_hd__buf_4
XFILLER_241_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26483_ _10798_ registers\[42\]\[32\] _11547_ VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23695_ _10011_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28222_ _11847_ registers\[30\]\[56\] _12490_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__mux2_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25434_ _10838_ registers\[50\]\[51\] _10992_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__mux2_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22646_ registers\[52\]\[56\] registers\[53\]\[56\] registers\[54\]\[56\] registers\[55\]\[56\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__mux4_1
XFILLER_224_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1053 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28153_ _11778_ registers\[30\]\[23\] _12457_ VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__mux2_1
X_25365_ _10957_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__clkbuf_1
X_22577_ _09218_ _09221_ _09083_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27104_ _11811_ registers\[38\]\[39\] _11898_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__mux2_1
X_24316_ _10352_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
X_28084_ _12424_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__clkbuf_1
X_21528_ registers\[8\]\[24\] registers\[9\]\[24\] registers\[10\]\[24\] registers\[11\]\[24\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__mux4_1
X_25296_ _10835_ registers\[51\]\[50\] _10920_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__mux2_1
XFILLER_166_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27035_ _11742_ registers\[38\]\[6\] _11865_ VGND VGND VPWR VPWR _11872_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24247_ registers\[57\]\[0\] _10303_ _10305_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__mux2_1
X_21459_ registers\[52\]\[22\] registers\[53\]\[22\] registers\[54\]\[22\] registers\[55\]\[22\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__mux4_1
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24178_ _09582_ registers\[58\]\[32\] _10266_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__mux2_1
XTAP_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23129_ _09686_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
XTAP_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28986_ registers\[24\]\[34\] _10376_ _12894_ VGND VGND VPWR VPWR _12899_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_62__f_CLK clknet_5_31_0_CLK VGND VGND VPWR VPWR clknet_6_62__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput97 net97 VGND VGND VPWR VPWR D1[16] sky130_fd_sc_hd__buf_2
XTAP_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27937_ registers\[32\]\[49\] _10407_ _12337_ VGND VGND VPWR VPWR _12347_ sky130_fd_sc_hd__mux2_1
XFILLER_7_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18670_ registers\[4\]\[8\] registers\[5\]\[8\] registers\[6\]\[8\] registers\[7\]\[8\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux4_1
XTAP_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27868_ registers\[32\]\[16\] _10338_ _12304_ VGND VGND VPWR VPWR _12311_ sky130_fd_sc_hd__mux2_1
XTAP_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ registers\[44\]\[44\] registers\[45\]\[44\] registers\[46\]\[44\] registers\[47\]\[44\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__mux4_1
X_29607_ registers\[20\]\[41\] _13021_ _13255_ VGND VGND VPWR VPWR _13257_ sky130_fd_sc_hd__mux2_1
XFILLER_40_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26819_ registers\[40\]\[63\] _10436_ _11657_ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__mux2_1
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27799_ _12274_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__clkbuf_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_406_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_406_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29538_ _13220_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__clkbuf_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ registers\[32\]\[42\] registers\[33\]\[42\] registers\[34\]\[42\] registers\[35\]\[42\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__mux4_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_940 _10303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_951 _10428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16503_ registers\[48\]\[12\] registers\[49\]\[12\] registers\[50\]\[12\] registers\[51\]\[12\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15005_ sky130_fd_sc_hd__mux4_1
XANTENNA_962 _10852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17483_ registers\[56\]\[40\] registers\[57\]\[40\] registers\[58\]\[40\] registers\[59\]\[40\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _15957_ sky130_fd_sc_hd__mux4_1
XFILLER_229_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29469_ _13139_ VGND VGND VPWR VPWR _13184_ sky130_fd_sc_hd__buf_4
XFILLER_225_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_973 _11158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_984 _11371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_31500_ _09780_ registers\[6\]\[42\] _14250_ VGND VGND VPWR VPWR _14253_ sky130_fd_sc_hd__mux2_1
XANTENNA_995 _11792_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19222_ _05747_ _05959_ _05960_ _05753_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a22o_1
X_16434_ _14562_ VGND VGND VPWR VPWR _14938_ sky130_fd_sc_hd__buf_6
XFILLER_38_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32480_ clknet_leaf_444_CLK _00594_ VGND VGND VPWR VPWR registers\[60\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16365_ registers\[0\]\[8\] registers\[1\]\[8\] registers\[2\]\[8\] registers\[3\]\[8\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14871_ sky130_fd_sc_hd__mux4_1
X_31431_ _14216_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__clkbuf_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19153_ _05890_ _05891_ _05892_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__a22o_1
XFILLER_188_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18104_ _14587_ _04871_ _04872_ _14597_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a22o_1
XFILLER_173_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34150_ clknet_leaf_432_CLK _02264_ VGND VGND VPWR VPWR registers\[34\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31362_ _14180_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__clkbuf_1
X_16296_ _14581_ VGND VGND VPWR VPWR _14804_ sky130_fd_sc_hd__buf_4
X_19084_ _05104_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__clkbuf_4
X_30313_ registers\[15\]\[56\] _13052_ _13621_ VGND VGND VPWR VPWR _13628_ sky130_fd_sc_hd__mux2_1
X_33101_ clknet_leaf_170_CLK _01215_ VGND VGND VPWR VPWR registers\[51\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_18035_ registers\[40\]\[56\] registers\[41\]\[56\] registers\[42\]\[56\] registers\[43\]\[56\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__mux4_1
XFILLER_172_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31293_ registers\[7\]\[8\] net63 _14135_ VGND VGND VPWR VPWR _14144_ sky130_fd_sc_hd__mux2_1
X_34081_ clknet_leaf_41_CLK _02195_ VGND VGND VPWR VPWR registers\[35\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33032_ clknet_leaf_192_CLK _01146_ VGND VGND VPWR VPWR registers\[52\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_30244_ registers\[15\]\[23\] _12983_ _13588_ VGND VGND VPWR VPWR _13592_ sky130_fd_sc_hd__mux2_1
XFILLER_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30175_ _13555_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__clkbuf_1
X_19986_ _06569_ _06701_ _06702_ _06574_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__a22o_1
XFILLER_154_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _05097_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__buf_4
X_34983_ clknet_leaf_457_CLK _03097_ VGND VGND VPWR VPWR registers\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1350 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1361 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1372 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33934_ clknet_leaf_132_CLK _02048_ VGND VGND VPWR VPWR registers\[37\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1383 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18868_ registers\[48\]\[14\] registers\[49\]\[14\] registers\[50\]\[14\] registers\[51\]\[14\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__mux4_1
XANTENNA_1394 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17819_ _04289_ _04595_ _04596_ _04292_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__a22o_1
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33865_ clknet_leaf_218_CLK _01979_ VGND VGND VPWR VPWR registers\[3\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_18799_ _05130_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__clkbuf_4
X_35604_ clknet_leaf_80_CLK _03718_ VGND VGND VPWR VPWR registers\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32816_ clknet_leaf_368_CLK _00930_ VGND VGND VPWR VPWR registers\[55\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_20830_ _07349_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__buf_4
X_33796_ clknet_leaf_252_CLK _01910_ VGND VGND VPWR VPWR registers\[40\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35535_ clknet_leaf_138_CLK _03649_ VGND VGND VPWR VPWR registers\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20761_ _07355_ _07456_ _07457_ _07367_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__a22o_1
X_32747_ clknet_leaf_420_CLK _00861_ VGND VGND VPWR VPWR registers\[56\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22500_ _09147_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35466_ clknet_leaf_150_CLK _03580_ VGND VGND VPWR VPWR registers\[14\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_23480_ _09567_ registers\[19\]\[25\] _09892_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__mux2_1
XFILLER_91_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20692_ _07315_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__buf_4
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32678_ clknet_leaf_439_CLK _00792_ VGND VGND VPWR VPWR registers\[57\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22431_ registers\[44\]\[50\] registers\[45\]\[50\] registers\[46\]\[50\] registers\[47\]\[50\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__mux4_1
X_34417_ clknet_leaf_386_CLK _02531_ VGND VGND VPWR VPWR registers\[30\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_31629_ _14320_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__clkbuf_1
X_35397_ clknet_leaf_228_CLK _03511_ VGND VGND VPWR VPWR registers\[15\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25150_ net47 VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__buf_2
XFILLER_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22362_ _07316_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__clkbuf_4
X_34348_ clknet_leaf_403_CLK _02462_ VGND VGND VPWR VPWR registers\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_248_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24101_ _10227_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21313_ registers\[52\]\[18\] registers\[53\]\[18\] registers\[54\]\[18\] registers\[55\]\[18\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__mux4_1
X_25081_ net22 VGND VGND VPWR VPWR _10791_ sky130_fd_sc_hd__buf_2
X_22293_ _08669_ _08944_ _08945_ _08675_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a22o_1
X_34279_ clknet_leaf_430_CLK _02393_ VGND VGND VPWR VPWR registers\[32\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24032_ _10191_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__clkbuf_1
X_36018_ clknet_leaf_380_CLK _04132_ VGND VGND VPWR VPWR registers\[63\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21244_ _07352_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__buf_4
XFILLER_11_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28840_ _11790_ registers\[25\]\[29\] _12812_ VGND VGND VPWR VPWR _12822_ sky130_fd_sc_hd__mux2_1
X_21175_ registers\[8\]\[14\] registers\[9\]\[14\] registers\[10\]\[14\] registers\[11\]\[14\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__mux4_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20126_ registers\[40\]\[50\] registers\[41\]\[50\] registers\[42\]\[50\] registers\[43\]\[50\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28771_ _12785_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25983_ _10838_ registers\[46\]\[51\] _11285_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__mux2_1
XFILLER_120_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20057_ registers\[44\]\[48\] registers\[45\]\[48\] registers\[46\]\[48\] registers\[47\]\[48\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__mux4_1
X_27722_ _12234_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__clkbuf_1
X_24934_ _10699_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24865_ _10663_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
X_27653_ registers\[34\]\[42\] _10393_ _12195_ VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__mux2_1
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23816_ _09628_ registers\[29\]\[54\] _10072_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__mux2_1
X_26604_ _10783_ registers\[41\]\[25\] _11608_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__mux2_1
XANTENNA_203 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27584_ _12161_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_214 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24796_ _09590_ registers\[54\]\[36\] _10620_ VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__mux2_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_236 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26535_ _10850_ registers\[42\]\[57\] _11569_ VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__mux2_1
XANTENNA_247 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29323_ _13107_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__clkbuf_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23747_ _09559_ registers\[29\]\[21\] _10039_ VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__mux2_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20959_ registers\[60\]\[8\] registers\[61\]\[8\] registers\[62\]\[8\] registers\[63\]\[8\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__mux4_1
XFILLER_42_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29254_ _13071_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__clkbuf_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26466_ _10781_ registers\[42\]\[24\] _11536_ VGND VGND VPWR VPWR _11541_ sky130_fd_sc_hd__mux2_1
X_23678_ registers\[61\]\[54\] _09806_ _09998_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__mux2_1
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28205_ _11830_ registers\[30\]\[48\] _12479_ VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__mux2_1
X_25417_ _10821_ registers\[50\]\[43\] _10981_ VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__mux2_1
X_22629_ registers\[28\]\[55\] registers\[29\]\[55\] registers\[30\]\[55\] registers\[31\]\[55\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__mux4_1
X_29185_ net38 VGND VGND VPWR VPWR _13025_ sky130_fd_sc_hd__buf_2
X_26397_ _11504_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16150_ registers\[48\]\[2\] registers\[49\]\[2\] registers\[50\]\[2\] registers\[51\]\[2\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14662_ sky130_fd_sc_hd__mux4_1
XFILLER_155_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28136_ _11761_ registers\[30\]\[15\] _12446_ VGND VGND VPWR VPWR _12452_ sky130_fd_sc_hd__mux2_1
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25348_ _10751_ registers\[50\]\[10\] _10948_ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__mux2_1
XFILLER_195_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16081_ _14594_ VGND VGND VPWR VPWR _14595_ sky130_fd_sc_hd__buf_4
X_28067_ _12415_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__clkbuf_1
X_25279_ _10819_ registers\[51\]\[42\] _10909_ VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__mux2_1
XFILLER_155_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27018_ _11861_ registers\[3\]\[63\] _11729_ VGND VGND VPWR VPWR _11862_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19840_ registers\[16\]\[41\] registers\[17\]\[41\] registers\[18\]\[41\] registers\[19\]\[41\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__mux4_1
XFILLER_155_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19771_ _06473_ _06480_ _06487_ _06494_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__or4_2
XFILLER_231_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28969_ registers\[24\]\[26\] _10359_ _12883_ VGND VGND VPWR VPWR _12890_ sky130_fd_sc_hd__mux2_1
X_16983_ _15341_ _15469_ _15470_ _15344_ VGND VGND VPWR VPWR _15471_ sky130_fd_sc_hd__a22o_1
XFILLER_231_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18722_ _05073_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__clkbuf_4
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31980_ clknet_leaf_4_CLK _00151_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18653_ _05045_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30931_ _13953_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__clkbuf_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17604_ _14520_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__buf_4
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33650_ clknet_leaf_360_CLK _01764_ VGND VGND VPWR VPWR registers\[42\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_30862_ _09819_ registers\[11\]\[60\] _13850_ VGND VGND VPWR VPWR _13917_ sky130_fd_sc_hd__mux2_1
XFILLER_184_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18584_ _05097_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__clkbuf_4
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32601_ clknet_leaf_84_CLK _00715_ VGND VGND VPWR VPWR registers\[58\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17535_ registers\[12\]\[41\] registers\[13\]\[41\] registers\[14\]\[41\] registers\[15\]\[41\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__mux4_1
X_33581_ clknet_leaf_318_CLK _01695_ VGND VGND VPWR VPWR registers\[43\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_30793_ _09747_ registers\[11\]\[27\] _13873_ VGND VGND VPWR VPWR _13881_ sky130_fd_sc_hd__mux2_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_770 _07835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35320_ clknet_leaf_309_CLK _03434_ VGND VGND VPWR VPWR registers\[16\]\[42\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_781 _08512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32532_ clknet_leaf_82_CLK _00646_ VGND VGND VPWR VPWR registers\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_792 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17466_ _15633_ _15939_ _15940_ _15636_ VGND VGND VPWR VPWR _15941_ sky130_fd_sc_hd__a22o_1
XFILLER_34_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19205_ _05839_ _05943_ _05944_ _05842_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__a22o_1
XFILLER_60_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16417_ _14502_ VGND VGND VPWR VPWR _14921_ sky130_fd_sc_hd__buf_4
X_35251_ clknet_leaf_409_CLK _03365_ VGND VGND VPWR VPWR registers\[17\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_32463_ clknet_leaf_175_CLK _00577_ VGND VGND VPWR VPWR registers\[60\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17397_ _15638_ _15872_ _15873_ _15643_ VGND VGND VPWR VPWR _15874_ sky130_fd_sc_hd__a22o_1
X_34202_ clknet_leaf_18_CLK _02316_ VGND VGND VPWR VPWR registers\[33\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_31414_ _09660_ registers\[6\]\[1\] _14206_ VGND VGND VPWR VPWR _14208_ sky130_fd_sc_hd__mux2_1
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19136_ registers\[28\]\[21\] registers\[29\]\[21\] registers\[30\]\[21\] registers\[31\]\[21\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__mux4_1
X_16348_ _14850_ _14853_ _14525_ VGND VGND VPWR VPWR _14854_ sky130_fd_sc_hd__o21ba_2
XFILLER_203_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35182_ clknet_leaf_397_CLK _03296_ VGND VGND VPWR VPWR registers\[18\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_32394_ clknet_leaf_177_CLK _00508_ VGND VGND VPWR VPWR registers\[61\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34133_ clknet_leaf_121_CLK _02247_ VGND VGND VPWR VPWR registers\[34\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16279_ registers\[56\]\[6\] registers\[57\]\[6\] registers\[58\]\[6\] registers\[59\]\[6\]
+ _14723_ _14532_ VGND VGND VPWR VPWR _14787_ sky130_fd_sc_hd__mux4_1
XFILLER_12_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31345_ _14171_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__clkbuf_1
X_19067_ registers\[40\]\[20\] registers\[41\]\[20\] registers\[42\]\[20\] registers\[43\]\[20\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__mux4_1
XFILLER_161_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18018_ _04786_ _04789_ _04619_ _04620_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__o211a_1
X_34064_ clknet_leaf_127_CLK _02178_ VGND VGND VPWR VPWR registers\[35\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31276_ _14134_ VGND VGND VPWR VPWR _14135_ sky130_fd_sc_hd__buf_4
X_33015_ clknet_leaf_328_CLK _01129_ VGND VGND VPWR VPWR registers\[52\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_30227_ registers\[15\]\[15\] _12966_ _13577_ VGND VGND VPWR VPWR _13583_ sky130_fd_sc_hd__mux2_1
XFILLER_82_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30158_ _13546_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19969_ registers\[0\]\[45\] registers\[1\]\[45\] registers\[2\]\[45\] registers\[3\]\[45\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__mux4_1
XFILLER_228_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34966_ clknet_leaf_97_CLK _03080_ VGND VGND VPWR VPWR registers\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_22980_ _09582_ registers\[62\]\[32\] _09578_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30089_ _13510_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1180 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1191 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33917_ clknet_leaf_276_CLK _02031_ VGND VGND VPWR VPWR registers\[38\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_21931_ registers\[40\]\[36\] registers\[41\]\[36\] registers\[42\]\[36\] registers\[43\]\[36\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__mux4_1
X_34897_ clknet_leaf_114_CLK _03011_ VGND VGND VPWR VPWR registers\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24650_ _10549_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33848_ clknet_leaf_316_CLK _01962_ VGND VGND VPWR VPWR registers\[3\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_21862_ _08524_ _08527_ _08430_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__o21ba_1
XFILLER_243_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23601_ _09962_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
X_20813_ _07314_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__buf_6
X_24581_ _10511_ VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__buf_12
X_21793_ _08439_ _08446_ _08453_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__or4_1
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33779_ clknet_leaf_346_CLK _01893_ VGND VGND VPWR VPWR registers\[40\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26320_ _10770_ registers\[43\]\[19\] _11454_ VGND VGND VPWR VPWR _11464_ sky130_fd_sc_hd__mux2_1
X_23532_ _09869_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__buf_4
XFILLER_196_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35518_ clknet_leaf_197_CLK _03632_ VGND VGND VPWR VPWR registers\[13\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_20744_ registers\[44\]\[2\] registers\[45\]\[2\] registers\[46\]\[2\] registers\[47\]\[2\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__mux4_1
XFILLER_223_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26251_ _10835_ registers\[44\]\[50\] _11427_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__mux2_1
X_35449_ clknet_leaf_304_CLK _03563_ VGND VGND VPWR VPWR registers\[14\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_23463_ _09550_ registers\[19\]\[17\] _09881_ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__mux2_1
X_20675_ _07361_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__buf_6
XFILLER_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25202_ _10871_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22414_ registers\[4\]\[49\] registers\[5\]\[49\] registers\[6\]\[49\] registers\[7\]\[49\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__mux4_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26182_ _11391_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
X_23394_ _09657_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__clkbuf_4
XFILLER_164_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25133_ _10826_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__clkbuf_1
X_22345_ registers\[24\]\[47\] registers\[25\]\[47\] registers\[26\]\[47\] registers\[27\]\[47\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__mux4_1
XFILLER_136_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29941_ _13432_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__clkbuf_1
X_25064_ _10779_ registers\[52\]\[23\] _10773_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__mux2_1
X_22276_ registers\[16\]\[45\] registers\[17\]\[45\] registers\[18\]\[45\] registers\[19\]\[45\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__mux4_1
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24015_ _10182_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21227_ _07776_ _07908_ _07909_ _07781_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__a22o_1
X_29872_ registers\[18\]\[39\] _13016_ _13386_ VGND VGND VPWR VPWR _13396_ sky130_fd_sc_hd__mux2_1
XFILLER_104_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28823_ _12813_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21158_ _07843_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20109_ _06819_ _06822_ _06512_ _06513_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__o211a_1
X_28754_ _11839_ registers\[26\]\[52\] _12774_ VGND VGND VPWR VPWR _12777_ sky130_fd_sc_hd__mux2_1
XFILLER_219_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25966_ _10821_ registers\[46\]\[43\] _11274_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__mux2_1
XFILLER_120_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21089_ _07312_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27705_ _12225_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24917_ _10690_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_833 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25897_ _10751_ registers\[46\]\[10\] _11241_ VGND VGND VPWR VPWR _11242_ sky130_fd_sc_hd__mux2_1
X_28685_ _12740_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__clkbuf_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27636_ registers\[34\]\[34\] _10376_ _12184_ VGND VGND VPWR VPWR _12189_ sky130_fd_sc_hd__mux2_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _09642_ registers\[54\]\[61\] _10586_ VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__mux2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27567_ registers\[34\]\[1\] _10307_ _12151_ VGND VGND VPWR VPWR _12153_ sky130_fd_sc_hd__mux2_1
XFILLER_26_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _09573_ registers\[54\]\[28\] _10609_ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__mux2_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17320_ _15487_ _15797_ _15798_ _15490_ VGND VGND VPWR VPWR _15799_ sky130_fd_sc_hd__a22o_1
X_29306_ _13098_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__clkbuf_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26518_ _10833_ registers\[42\]\[49\] _11558_ VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__mux2_1
XFILLER_18_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27498_ _12115_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29237_ net57 VGND VGND VPWR VPWR _13060_ sky130_fd_sc_hd__buf_2
XFILLER_186_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17251_ _14520_ VGND VGND VPWR VPWR _15732_ sky130_fd_sc_hd__buf_4
X_26449_ _10764_ registers\[42\]\[16\] _11525_ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__mux2_1
XFILLER_202_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16202_ _14601_ _14711_ _14712_ _14611_ VGND VGND VPWR VPWR _14713_ sky130_fd_sc_hd__a22o_1
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17182_ registers\[12\]\[31\] registers\[13\]\[31\] registers\[14\]\[31\] registers\[15\]\[31\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15665_ sky130_fd_sc_hd__mux4_1
XFILLER_35_1374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29168_ _13013_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16133_ _14642_ _14645_ _14614_ VGND VGND VPWR VPWR _14646_ sky130_fd_sc_hd__o21ba_1
X_28119_ _11744_ registers\[30\]\[7\] _12435_ VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__mux2_1
XFILLER_6_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29099_ registers\[23\]\[15\] _12966_ _12956_ VGND VGND VPWR VPWR _12967_ sky130_fd_sc_hd__mux2_1
XFILLER_170_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31130_ registers\[0\]\[59\] _13058_ _14048_ VGND VGND VPWR VPWR _14058_ sky130_fd_sc_hd__mux2_1
XFILLER_142_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16064_ _14531_ VGND VGND VPWR VPWR _14578_ sky130_fd_sc_hd__buf_12
XFILLER_192_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31061_ registers\[0\]\[26\] _12989_ _14015_ VGND VGND VPWR VPWR _14022_ sky130_fd_sc_hd__mux2_1
XFILLER_123_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30012_ registers\[17\]\[41\] _13021_ _13468_ VGND VGND VPWR VPWR _13470_ sky130_fd_sc_hd__mux2_1
XFILLER_97_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19823_ _06233_ _06543_ _06544_ _06236_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__a22o_1
XFILLER_151_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34820_ clknet_leaf_225_CLK _02934_ VGND VGND VPWR VPWR registers\[24\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19754_ registers\[52\]\[39\] registers\[53\]\[39\] registers\[54\]\[39\] registers\[55\]\[39\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__mux4_1
X_16966_ registers\[4\]\[25\] registers\[5\]\[25\] registers\[6\]\[25\] registers\[7\]\[25\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15455_ sky130_fd_sc_hd__mux4_1
XFILLER_231_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18705_ registers\[24\]\[9\] registers\[25\]\[9\] registers\[26\]\[9\] registers\[27\]\[9\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__mux4_1
X_34751_ clknet_leaf_189_CLK _02865_ VGND VGND VPWR VPWR registers\[25\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_31963_ clknet_leaf_4_CLK _00132_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
X_19685_ registers\[8\]\[37\] registers\[9\]\[37\] registers\[10\]\[37\] registers\[11\]\[37\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__mux4_1
X_16897_ _14518_ VGND VGND VPWR VPWR _15388_ sky130_fd_sc_hd__buf_4
X_33702_ clknet_leaf_430_CLK _01816_ VGND VGND VPWR VPWR registers\[41\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18636_ registers\[28\]\[7\] registers\[29\]\[7\] registers\[30\]\[7\] registers\[31\]\[7\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__mux4_1
X_30914_ registers\[10\]\[20\] _12976_ _13944_ VGND VGND VPWR VPWR _13945_ sky130_fd_sc_hd__mux2_1
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34682_ clknet_leaf_184_CLK _02796_ VGND VGND VPWR VPWR registers\[26\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31894_ _09769_ registers\[49\]\[37\] _14452_ VGND VGND VPWR VPWR _14460_ sky130_fd_sc_hd__mux2_1
XFILLER_224_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33633_ clknet_leaf_33_CLK _01747_ VGND VGND VPWR VPWR registers\[42\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_30845_ _13908_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__clkbuf_1
X_18567_ registers\[20\]\[5\] registers\[21\]\[5\] registers\[22\]\[5\] registers\[23\]\[5\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__mux4_1
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17518_ registers\[40\]\[41\] registers\[41\]\[41\] registers\[42\]\[41\] registers\[43\]\[41\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__mux4_1
X_33564_ clknet_leaf_28_CLK _01678_ VGND VGND VPWR VPWR registers\[43\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18498_ registers\[16\]\[3\] registers\[17\]\[3\] registers\[18\]\[3\] registers\[19\]\[3\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__mux4_1
X_30776_ _09697_ registers\[11\]\[19\] _13862_ VGND VGND VPWR VPWR _13872_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35303_ clknet_leaf_448_CLK _03417_ VGND VGND VPWR VPWR registers\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_32515_ clknet_leaf_293_CLK _00629_ VGND VGND VPWR VPWR registers\[60\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_17449_ _15920_ _15923_ _15612_ VGND VGND VPWR VPWR _15924_ sky130_fd_sc_hd__o21ba_1
X_33495_ clknet_leaf_123_CLK _01609_ VGND VGND VPWR VPWR registers\[44\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35234_ clknet_leaf_474_CLK _03348_ VGND VGND VPWR VPWR registers\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_20460_ _06919_ _07161_ _07162_ _06922_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__a22o_1
X_32446_ clknet_leaf_183_CLK _00560_ VGND VGND VPWR VPWR registers\[29\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19119_ registers\[56\]\[21\] registers\[57\]\[21\] registers\[58\]\[21\] registers\[59\]\[21\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__mux4_1
X_35165_ clknet_leaf_5_CLK _03279_ VGND VGND VPWR VPWR registers\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20391_ _06873_ _07095_ _07096_ _06878_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__a22o_1
XFILLER_174_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32377_ clknet_leaf_332_CLK _00491_ VGND VGND VPWR VPWR registers\[61\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34116_ clknet_leaf_246_CLK _02230_ VGND VGND VPWR VPWR registers\[35\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_22130_ _08677_ _08786_ _08787_ _08681_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__a22o_1
X_31328_ _14162_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput210 net210 VGND VGND VPWR VPWR D2[60] sky130_fd_sc_hd__buf_2
X_35096_ clknet_leaf_11_CLK _03210_ VGND VGND VPWR VPWR registers\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xoutput221 net221 VGND VGND VPWR VPWR D3[12] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR D3[22] sky130_fd_sc_hd__buf_2
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34047_ clknet_leaf_275_CLK _02161_ VGND VGND VPWR VPWR registers\[36\]\[49\] sky130_fd_sc_hd__dfxtp_1
Xoutput243 net243 VGND VGND VPWR VPWR D3[32] sky130_fd_sc_hd__buf_2
X_22061_ registers\[4\]\[39\] registers\[5\]\[39\] registers\[6\]\[39\] registers\[7\]\[39\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__mux4_1
XTAP_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31259_ registers\[8\]\[56\] net52 _14119_ VGND VGND VPWR VPWR _14126_ sky130_fd_sc_hd__mux2_1
Xoutput254 net254 VGND VGND VPWR VPWR D3[42] sky130_fd_sc_hd__buf_2
XFILLER_82_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput265 net265 VGND VGND VPWR VPWR D3[52] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR D3[62] sky130_fd_sc_hd__buf_2
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21012_ _07680_ _07687_ _07694_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__or4_1
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25820_ _10810_ registers\[47\]\[38\] _11192_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__mux2_1
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35998_ clknet_leaf_46_CLK _04112_ VGND VGND VPWR VPWR registers\[63\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25751_ _10741_ registers\[47\]\[5\] _11159_ VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34949_ clknet_leaf_205_CLK _03063_ VGND VGND VPWR VPWR registers\[22\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_22963_ net20 VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__buf_2
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24702_ _10576_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
X_21914_ _07289_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__buf_4
XFILLER_215_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28470_ _12627_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__clkbuf_1
X_25682_ _11127_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
X_22894_ _09524_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27421_ _12074_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24633_ _10540_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
X_21845_ _08334_ _08509_ _08510_ _08338_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__a22o_1
XFILLER_231_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24564_ _10502_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27352_ _12038_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__clkbuf_1
X_21776_ registers\[52\]\[31\] registers\[53\]\[31\] registers\[54\]\[31\] registers\[55\]\[31\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__mux4_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26303_ _11455_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
X_23515_ _09916_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27283_ _11855_ registers\[37\]\[60\] _11935_ VGND VGND VPWR VPWR _12002_ sky130_fd_sc_hd__mux2_1
X_20727_ registers\[24\]\[1\] registers\[25\]\[1\] registers\[26\]\[1\] registers\[27\]\[1\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__mux4_1
X_24495_ _10466_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29022_ registers\[24\]\[51\] _10412_ _12916_ VGND VGND VPWR VPWR _12918_ sky130_fd_sc_hd__mux2_1
XFILLER_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26234_ _10819_ registers\[44\]\[42\] _11416_ VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__mux2_1
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23446_ _09533_ registers\[19\]\[9\] _09870_ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__mux2_1
X_20658_ _07356_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__buf_8
XFILLER_109_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26165_ _11382_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23377_ _09842_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
X_20589_ _07287_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__buf_4
XFILLER_165_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25116_ _10730_ VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__buf_4
X_22328_ registers\[36\]\[47\] registers\[37\]\[47\] registers\[38\]\[47\] registers\[39\]\[47\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__mux4_1
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26096_ _11346_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
X_29924_ _09707_ _12933_ VGND VGND VPWR VPWR _13423_ sky130_fd_sc_hd__nor2_8
X_25047_ net10 VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__clkbuf_4
X_22259_ registers\[56\]\[45\] registers\[57\]\[45\] registers\[58\]\[45\] registers\[59\]\[45\]
+ _08880_ _08670_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__mux4_1
XFILLER_219_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29855_ _13387_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28806_ _12804_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16820_ registers\[48\]\[21\] registers\[49\]\[21\] registers\[50\]\[21\] registers\[51\]\[21\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15313_ sky130_fd_sc_hd__mux4_1
X_29786_ _13350_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26998_ _11848_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28737_ _11822_ registers\[26\]\[44\] _12763_ VGND VGND VPWR VPWR _12768_ sky130_fd_sc_hd__mux2_1
X_16751_ registers\[8\]\[19\] registers\[9\]\[19\] registers\[10\]\[19\] registers\[11\]\[19\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15246_ sky130_fd_sc_hd__mux4_1
XFILLER_65_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25949_ _10804_ registers\[46\]\[35\] _11263_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19470_ _05890_ _06200_ _06201_ _05893_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__a22o_1
X_16682_ registers\[12\]\[17\] registers\[13\]\[17\] registers\[14\]\[17\] registers\[15\]\[17\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15179_ sky130_fd_sc_hd__mux4_1
X_28668_ _11753_ registers\[26\]\[11\] _12730_ VGND VGND VPWR VPWR _12732_ sky130_fd_sc_hd__mux2_1
X_18421_ registers\[0\]\[1\] registers\[1\]\[1\] registers\[2\]\[1\] registers\[3\]\[1\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__mux4_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27619_ registers\[34\]\[26\] _10359_ _12173_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28599_ _12695_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ registers\[0\]\[0\] registers\[1\]\[0\] registers\[2\]\[0\] registers\[3\]\[0\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__mux4_1
X_30630_ _13795_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__clkbuf_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ registers\[36\]\[35\] registers\[37\]\[35\] registers\[38\]\[35\] registers\[39\]\[35\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15782_ sky130_fd_sc_hd__mux4_1
XFILLER_230_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18283_ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__clkbuf_8
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30561_ _09786_ registers\[13\]\[45\] _13753_ VGND VGND VPWR VPWR _13759_ sky130_fd_sc_hd__mux2_1
XFILLER_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32300_ clknet_leaf_396_CLK _00414_ VGND VGND VPWR VPWR registers\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_17234_ registers\[32\]\[33\] registers\[33\]\[33\] registers\[34\]\[33\] registers\[35\]\[33\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15715_ sky130_fd_sc_hd__mux4_1
X_33280_ clknet_leaf_270_CLK _01394_ VGND VGND VPWR VPWR registers\[48\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30492_ _09683_ registers\[13\]\[12\] _13720_ VGND VGND VPWR VPWR _13723_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32231_ clknet_leaf_151_CLK _00345_ VGND VGND VPWR VPWR registers\[9\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17165_ registers\[40\]\[31\] registers\[41\]\[31\] registers\[42\]\[31\] registers\[43\]\[31\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15648_ sky130_fd_sc_hd__mux4_1
X_16116_ registers\[60\]\[1\] registers\[61\]\[1\] registers\[62\]\[1\] registers\[63\]\[1\]
+ _14542_ _14544_ VGND VGND VPWR VPWR _14629_ sky130_fd_sc_hd__mux4_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32162_ clknet_leaf_440_CLK _00276_ VGND VGND VPWR VPWR registers\[39\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17096_ _15577_ _15580_ _15269_ VGND VGND VPWR VPWR _15581_ sky130_fd_sc_hd__o21ba_1
XFILLER_182_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31113_ _14049_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16047_ registers\[8\]\[0\] registers\[9\]\[0\] registers\[10\]\[0\] registers\[11\]\[0\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _14561_ sky130_fd_sc_hd__mux4_1
X_32093_ clknet_leaf_485_CLK _00006_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35921_ clknet_leaf_107_CLK _04035_ VGND VGND VPWR VPWR registers\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31044_ registers\[0\]\[18\] _12972_ _14004_ VGND VGND VPWR VPWR _14013_ sky130_fd_sc_hd__mux2_1
XFILLER_215_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19806_ _06525_ _06526_ _06527_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__a22o_1
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35852_ clknet_leaf_144_CLK _03966_ VGND VGND VPWR VPWR registers\[8\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17998_ _04632_ _04769_ _04770_ _04635_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__a22o_1
XFILLER_215_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34803_ clknet_leaf_414_CLK _02917_ VGND VGND VPWR VPWR registers\[24\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_19737_ _06187_ _06460_ _06461_ _06192_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__a22o_1
X_35783_ clknet_leaf_217_CLK _03897_ VGND VGND VPWR VPWR registers\[0\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_16949_ registers\[44\]\[25\] registers\[45\]\[25\] registers\[46\]\[25\] registers\[47\]\[25\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15438_ sky130_fd_sc_hd__mux4_1
X_32995_ clknet_leaf_441_CLK _01109_ VGND VGND VPWR VPWR registers\[52\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_34734_ clknet_leaf_411_CLK _02848_ VGND VGND VPWR VPWR registers\[25\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_31946_ _09823_ registers\[49\]\[62\] _14418_ VGND VGND VPWR VPWR _14487_ sky130_fd_sc_hd__mux2_1
X_19668_ _06394_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__buf_2
XFILLER_225_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18619_ registers\[56\]\[7\] registers\[57\]\[7\] registers\[58\]\[7\] registers\[59\]\[7\]
+ _05272_ _05081_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__mux4_1
XFILLER_213_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34665_ clknet_leaf_452_CLK _02779_ VGND VGND VPWR VPWR registers\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_19599_ registers\[40\]\[35\] registers\[41\]\[35\] registers\[42\]\[35\] registers\[43\]\[35\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__mux4_1
X_31877_ _09751_ registers\[49\]\[29\] _14441_ VGND VGND VPWR VPWR _14451_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33616_ clknet_leaf_128_CLK _01730_ VGND VGND VPWR VPWR registers\[42\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_39__f_CLK clknet_5_19_0_CLK VGND VGND VPWR VPWR clknet_6_39__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_21630_ _07991_ _08300_ _08301_ _07995_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__a22o_1
X_30828_ _13899_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__clkbuf_1
X_34596_ clknet_leaf_445_CLK _02710_ VGND VGND VPWR VPWR registers\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33547_ clknet_leaf_163_CLK _01661_ VGND VGND VPWR VPWR registers\[44\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21561_ _07289_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__buf_4
X_30759_ _13863_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23300_ net44 VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__clkbuf_4
X_20512_ _07210_ _07213_ _05162_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__o21ba_1
X_24280_ net3 VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__buf_4
X_33478_ clknet_leaf_254_CLK _01592_ VGND VGND VPWR VPWR registers\[45\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21492_ _07991_ _08166_ _08167_ _07995_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__a22o_1
X_35217_ clknet_leaf_113_CLK _03331_ VGND VGND VPWR VPWR registers\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_23231_ net21 VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__buf_4
X_20443_ registers\[4\]\[59\] registers\[5\]\[59\] registers\[6\]\[59\] registers\[7\]\[59\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__mux4_1
X_32429_ clknet_leaf_396_CLK _00543_ VGND VGND VPWR VPWR registers\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36197_ clknet_leaf_98_CLK _00079_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35148_ clknet_leaf_149_CLK _03262_ VGND VGND VPWR VPWR registers\[1\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_23162_ _09710_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__clkbuf_1
X_20374_ _06776_ _07078_ _07079_ _06782_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22113_ _08766_ _08767_ _08770_ _08771_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__a22o_1
XTAP_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35079_ clknet_leaf_206_CLK _03193_ VGND VGND VPWR VPWR registers\[20\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_27970_ _11728_ registers\[31\]\[0\] _12364_ VGND VGND VPWR VPWR _12365_ sky130_fd_sc_hd__mux2_1
X_23093_ net23 VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__buf_4
XTAP_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26921_ _11796_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22044_ registers\[32\]\[39\] registers\[33\]\[39\] registers\[34\]\[39\] registers\[35\]\[39\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__mux4_1
XTAP_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29640_ registers\[20\]\[57\] _13054_ _13266_ VGND VGND VPWR VPWR _13274_ sky130_fd_sc_hd__mux2_1
XTAP_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26852_ _11749_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_1
XTAP_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25803_ _11158_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__buf_4
X_29571_ registers\[20\]\[24\] _12985_ _13233_ VGND VGND VPWR VPWR _13238_ sky130_fd_sc_hd__mux2_1
XFILLER_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26783_ _11708_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__clkbuf_1
X_23995_ _10160_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__buf_4
XFILLER_235_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28522_ _11742_ registers\[27\]\[6\] _12648_ VGND VGND VPWR VPWR _12655_ sky130_fd_sc_hd__mux2_1
XFILLER_84_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25734_ _11154_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
X_22946_ _09559_ registers\[62\]\[21\] _09557_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28453_ _12618_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__clkbuf_1
X_22877_ net88 net87 net86 net89 VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__and4_2
XFILLER_216_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25665_ _11118_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27404_ registers\[36\]\[53\] _10416_ _12062_ VGND VGND VPWR VPWR _12066_ sky130_fd_sc_hd__mux2_1
X_24616_ _10531_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
X_21828_ registers\[20\]\[32\] registers\[21\]\[32\] registers\[22\]\[32\] registers\[23\]\[32\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__mux4_1
XFILLER_19_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25596_ _11080_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28384_ _12582_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24547_ _10493_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
X_27335_ registers\[36\]\[20\] _10346_ _12029_ VGND VGND VPWR VPWR _12030_ sky130_fd_sc_hd__mux2_1
X_21759_ _07395_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27266_ _11993_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__clkbuf_1
X_24478_ _10457_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29005_ registers\[24\]\[43\] _10395_ _12905_ VGND VGND VPWR VPWR _12909_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23429_ _09871_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26217_ _10802_ registers\[44\]\[34\] _11405_ VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__mux2_1
X_27197_ _11769_ registers\[37\]\[19\] _11947_ VGND VGND VPWR VPWR _11957_ sky130_fd_sc_hd__mux2_1
XFILLER_125_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26148_ _10733_ registers\[44\]\[1\] _11372_ VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__mux2_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26079_ _11337_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
X_18970_ _05547_ _05712_ _05715_ _05550_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__a22o_1
XFILLER_180_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ registers\[8\]\[52\] registers\[9\]\[52\] registers\[10\]\[52\] registers\[11\]\[52\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__mux4_1
X_29907_ _13414_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__clkbuf_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1702 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1713 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1724 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1735 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1746 _05059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ _04486_ _04627_ _04628_ _04489_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a22o_1
XANTENNA_1757 _07316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29838_ _13378_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__clkbuf_1
XTAP_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1768 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1779 _12006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16803_ _14530_ VGND VGND VPWR VPWR _15297_ sky130_fd_sc_hd__buf_4
X_29769_ registers\[1\]\[54\] _13048_ _13337_ VGND VGND VPWR VPWR _13342_ sky130_fd_sc_hd__mux2_1
X_17783_ _04486_ _04558_ _04561_ _04489_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__a22o_1
XFILLER_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31800_ _14410_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__clkbuf_1
X_19522_ registers\[24\]\[32\] registers\[25\]\[32\] registers\[26\]\[32\] registers\[27\]\[32\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__mux4_1
XFILLER_208_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16734_ _15229_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32780_ clknet_leaf_167_CLK _00894_ VGND VGND VPWR VPWR registers\[56\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19453_ _06182_ _06183_ _06184_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a22o_1
X_31731_ _14374_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__clkbuf_1
X_16665_ _14991_ _15160_ _15161_ _14996_ VGND VGND VPWR VPWR _15162_ sky130_fd_sc_hd__a22o_1
XFILLER_235_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18404_ registers\[40\]\[1\] registers\[41\]\[1\] registers\[42\]\[1\] registers\[43\]\[1\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__mux4_1
XFILLER_223_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34450_ clknet_leaf_105_CLK _02564_ VGND VGND VPWR VPWR registers\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_31662_ registers\[63\]\[55\] net51 _14332_ VGND VGND VPWR VPWR _14338_ sky130_fd_sc_hd__mux2_1
X_19384_ _05844_ _06117_ _06118_ _05849_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a22o_1
XFILLER_37_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16596_ registers\[44\]\[15\] registers\[45\]\[15\] registers\[46\]\[15\] registers\[47\]\[15\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15095_ sky130_fd_sc_hd__mux4_1
XFILLER_210_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33401_ clknet_leaf_280_CLK _01515_ VGND VGND VPWR VPWR registers\[46\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_18335_ _05097_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__clkbuf_4
X_30613_ _13786_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__clkbuf_1
X_34381_ clknet_leaf_141_CLK _02495_ VGND VGND VPWR VPWR registers\[31\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31593_ registers\[63\]\[22\] net15 _14299_ VGND VGND VPWR VPWR _14302_ sky130_fd_sc_hd__mux2_1
XFILLER_175_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36120_ clknet_leaf_53_CLK _04234_ VGND VGND VPWR VPWR registers\[49\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33332_ clknet_leaf_345_CLK _01446_ VGND VGND VPWR VPWR registers\[47\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_18266_ registers\[24\]\[63\] registers\[25\]\[63\] registers\[26\]\[63\] registers\[27\]\[63\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux4_1
X_30544_ _09769_ registers\[13\]\[37\] _13742_ VGND VGND VPWR VPWR _13750_ sky130_fd_sc_hd__mux2_1
XFILLER_198_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36051_ clknet_leaf_71_CLK _04165_ VGND VGND VPWR VPWR registers\[59\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17217_ _15482_ _15697_ _15698_ _15485_ VGND VGND VPWR VPWR _15699_ sky130_fd_sc_hd__a22o_1
X_33263_ clknet_leaf_364_CLK _01377_ VGND VGND VPWR VPWR registers\[48\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_18197_ _14600_ _04961_ _04962_ _14610_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__a22o_1
X_30475_ _09666_ registers\[13\]\[4\] _13709_ VGND VGND VPWR VPWR _13714_ sky130_fd_sc_hd__mux2_1
XFILLER_11_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35002_ clknet_leaf_308_CLK _03116_ VGND VGND VPWR VPWR registers\[21\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_32214_ clknet_leaf_288_CLK _00328_ VGND VGND VPWR VPWR registers\[9\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_17148_ _15627_ _15630_ _15631_ VGND VGND VPWR VPWR _15632_ sky130_fd_sc_hd__o21ba_1
XFILLER_239_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33194_ clknet_leaf_402_CLK _01308_ VGND VGND VPWR VPWR registers\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32145_ clknet_leaf_134_CLK _00259_ VGND VGND VPWR VPWR registers\[39\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17079_ registers\[24\]\[28\] registers\[25\]\[28\] registers\[26\]\[28\] registers\[27\]\[28\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15565_ sky130_fd_sc_hd__mux4_1
XFILLER_83_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32076_ clknet_leaf_167_CLK _00254_ VGND VGND VPWR VPWR registers\[62\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_20090_ _06530_ _06803_ _06804_ _06535_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__a22o_1
XFILLER_131_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35904_ clknet_leaf_234_CLK _04018_ VGND VGND VPWR VPWR registers\[7\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_31027_ _13992_ VGND VGND VPWR VPWR _14004_ sky130_fd_sc_hd__buf_4
XFILLER_83_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35835_ clknet_leaf_288_CLK _03949_ VGND VGND VPWR VPWR registers\[8\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22800_ registers\[0\]\[61\] registers\[1\]\[61\] registers\[2\]\[61\] registers\[3\]\[61\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__mux4_1
XFILLER_211_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23780_ _09592_ registers\[29\]\[37\] _10050_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__mux2_1
X_32978_ clknet_leaf_173_CLK _01092_ VGND VGND VPWR VPWR registers\[52\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_20992_ registers\[48\]\[9\] registers\[49\]\[9\] registers\[50\]\[9\] registers\[51\]\[9\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__mux4_1
X_35766_ clknet_leaf_331_CLK _03880_ VGND VGND VPWR VPWR registers\[0\]\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22731_ _09367_ _09370_ _09083_ VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__o21ba_2
X_31929_ _14478_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34717_ clknet_leaf_9_CLK _02831_ VGND VGND VPWR VPWR registers\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35697_ clknet_leaf_381_CLK _03811_ VGND VGND VPWR VPWR registers\[10\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25450_ _10854_ registers\[50\]\[59\] _10992_ VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22662_ _09301_ _09304_ _09116_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__o21ba_1
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34648_ clknet_leaf_18_CLK _02762_ VGND VGND VPWR VPWR registers\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24401_ _10304_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__buf_6
X_21613_ _08282_ _08285_ _08087_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__o21ba_1
XFILLER_179_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25381_ _10785_ registers\[50\]\[26\] _10959_ VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__mux2_1
X_22593_ _09234_ _09237_ _09102_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__o21ba_1
X_34579_ clknet_leaf_104_CLK _02693_ VGND VGND VPWR VPWR registers\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27120_ _11916_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__clkbuf_1
X_24332_ net21 VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__buf_4
XFILLER_142_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21544_ _08193_ _08202_ _08209_ _08218_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__or4_4
XFILLER_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27051_ _11880_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__clkbuf_1
X_24263_ _10316_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
X_21475_ registers\[20\]\[22\] registers\[21\]\[22\] registers\[22\]\[22\] registers\[23\]\[22\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__mux4_1
X_26002_ _11296_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23214_ _09738_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
X_20426_ registers\[32\]\[59\] registers\[33\]\[59\] registers\[34\]\[59\] registers\[35\]\[59\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__mux4_1
XFILLER_135_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24194_ _10232_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__buf_4
X_23145_ net11 VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__buf_4
X_20357_ registers\[16\]\[56\] registers\[17\]\[56\] registers\[18\]\[56\] registers\[19\]\[56\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__mux4_1
XFILLER_218_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27953_ _12355_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1009 _11853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23076_ _09647_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20288_ registers\[0\]\[54\] registers\[1\]\[54\] registers\[2\]\[54\] registers\[3\]\[54\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__mux4_1
XTAP_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26904_ _11784_ registers\[3\]\[26\] _11772_ VGND VGND VPWR VPWR _11785_ sky130_fd_sc_hd__mux2_1
X_22027_ _07361_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_130_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_130_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27884_ _12319_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29623_ registers\[20\]\[49\] _13037_ _13255_ VGND VGND VPWR VPWR _13265_ sky130_fd_sc_hd__mux2_1
XTAP_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26835_ net45 VGND VGND VPWR VPWR _11738_ sky130_fd_sc_hd__buf_4
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29554_ registers\[20\]\[16\] _12968_ _13222_ VGND VGND VPWR VPWR _13229_ sky130_fd_sc_hd__mux2_1
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26766_ _11699_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__clkbuf_1
X_23978_ _10163_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28505_ _12645_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25717_ registers\[48\]\[54\] _10418_ _11141_ VGND VGND VPWR VPWR _11146_ sky130_fd_sc_hd__mux2_1
X_29485_ _13192_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__clkbuf_1
X_22929_ net8 VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__buf_4
X_26697_ _11663_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28436_ _12609_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__clkbuf_1
X_16450_ _14530_ VGND VGND VPWR VPWR _14954_ sky130_fd_sc_hd__buf_4
XFILLER_204_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25648_ registers\[48\]\[21\] _10349_ _11108_ VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__mux2_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28367_ registers\[2\]\[61\] _10432_ _12505_ VGND VGND VPWR VPWR _12573_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_22__f_CLK clknet_5_11_0_CLK VGND VGND VPWR VPWR clknet_6_22__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_197_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_197_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16381_ _14886_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
X_25579_ registers\[4\]\[54\] _10418_ _11067_ VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__mux2_1
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18120_ registers\[20\]\[58\] registers\[21\]\[58\] registers\[22\]\[58\] registers\[23\]\[58\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__mux4_1
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27318_ registers\[36\]\[12\] _10330_ _12018_ VGND VGND VPWR VPWR _12021_ sky130_fd_sc_hd__mux2_1
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28298_ registers\[2\]\[28\] _10363_ _12528_ VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__mux2_1
XFILLER_40_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18051_ _14491_ _04820_ _04821_ _14501_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__a22o_1
XFILLER_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27249_ _11984_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17002_ _14581_ VGND VGND VPWR VPWR _15490_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30260_ _13600_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30191_ _13563_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18953_ _05141_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__buf_6
XFILLER_193_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1510 _07395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1521 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17904_ registers\[40\]\[52\] registers\[41\]\[52\] registers\[42\]\[52\] registers\[43\]\[52\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__mux4_1
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1532 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33950_ clknet_leaf_23_CLK _02064_ VGND VGND VPWR VPWR registers\[37\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_121_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_121_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_1543 _10232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18884_ registers\[24\]\[14\] registers\[25\]\[14\] registers\[26\]\[14\] registers\[27\]\[14\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__mux4_1
XTAP_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1554 _11513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1565 _11864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32901_ clknet_leaf_200_CLK _01015_ VGND VGND VPWR VPWR registers\[54\]\[55\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1576 _13637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17835_ _04605_ _04610_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1587 _14493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33881_ clknet_leaf_29_CLK _01995_ VGND VGND VPWR VPWR registers\[38\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1598 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32832_ clknet_leaf_294_CLK _00946_ VGND VGND VPWR VPWR registers\[55\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_35620_ clknet_leaf_465_CLK _03734_ VGND VGND VPWR VPWR registers\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17766_ registers\[48\]\[48\] registers\[49\]\[48\] registers\[50\]\[48\] registers\[51\]\[48\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__mux4_1
X_19505_ _05065_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_235_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35551_ clknet_leaf_482_CLK _03665_ VGND VGND VPWR VPWR registers\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16717_ registers\[8\]\[18\] registers\[9\]\[18\] registers\[10\]\[18\] registers\[11\]\[18\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15213_ sky130_fd_sc_hd__mux4_1
X_32763_ clknet_leaf_284_CLK _00877_ VGND VGND VPWR VPWR registers\[56\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17697_ registers\[52\]\[46\] registers\[53\]\[46\] registers\[54\]\[46\] registers\[55\]\[46\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__mux4_1
XFILLER_235_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34502_ clknet_leaf_217_CLK _02616_ VGND VGND VPWR VPWR registers\[2\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19436_ _05102_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__clkbuf_4
X_31714_ _14365_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__clkbuf_1
X_16648_ registers\[4\]\[16\] registers\[5\]\[16\] registers\[6\]\[16\] registers\[7\]\[16\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15146_ sky130_fd_sc_hd__mux4_1
X_35482_ clknet_leaf_13_CLK _03596_ VGND VGND VPWR VPWR registers\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32694_ clknet_leaf_334_CLK _00808_ VGND VGND VPWR VPWR registers\[57\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34433_ clknet_leaf_203_CLK _02547_ VGND VGND VPWR VPWR registers\[30\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_188_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_188_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31645_ registers\[63\]\[47\] net42 _14321_ VGND VGND VPWR VPWR _14329_ sky130_fd_sc_hd__mux2_1
X_19367_ _05065_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__buf_4
XFILLER_241_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16579_ registers\[4\]\[14\] registers\[5\]\[14\] registers\[6\]\[14\] registers\[7\]\[14\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15079_ sky130_fd_sc_hd__mux4_1
XFILLER_194_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18318_ _05080_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__buf_4
X_34364_ clknet_leaf_187_CLK _02478_ VGND VGND VPWR VPWR registers\[31\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31576_ registers\[63\]\[14\] net6 _14288_ VGND VGND VPWR VPWR _14293_ sky130_fd_sc_hd__mux2_1
X_19298_ _06031_ _06032_ _06033_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__a22o_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36103_ clknet_leaf_262_CLK _04217_ VGND VGND VPWR VPWR registers\[59\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33315_ clknet_leaf_57_CLK _01429_ VGND VGND VPWR VPWR registers\[47\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_18249_ registers\[36\]\[63\] registers\[37\]\[63\] registers\[38\]\[63\] registers\[39\]\[63\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__mux4_1
X_30527_ _09751_ registers\[13\]\[29\] _13731_ VGND VGND VPWR VPWR _13741_ sky130_fd_sc_hd__mux2_1
X_34295_ clknet_leaf_341_CLK _02409_ VGND VGND VPWR VPWR registers\[32\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36034_ clknet_leaf_264_CLK _04148_ VGND VGND VPWR VPWR registers\[63\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21260_ _07939_ _07942_ _07744_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__o21ba_1
XFILLER_89_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33246_ clknet_leaf_39_CLK _01360_ VGND VGND VPWR VPWR registers\[48\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30458_ _13704_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20211_ _05065_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__buf_4
XFILLER_239_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33177_ clknet_leaf_475_CLK _01291_ VGND VGND VPWR VPWR registers\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_360_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_360_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21191_ _07850_ _07859_ _07866_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__or4_2
XFILLER_144_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30389_ _13668_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20142_ _05102_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__clkbuf_4
X_32128_ clknet_leaf_397_CLK _00045_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dfxtp_1
XFILLER_132_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_112_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20073_ _05064_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__buf_4
X_32059_ clknet_leaf_287_CLK _00237_ VGND VGND VPWR VPWR registers\[62\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_24950_ _09609_ registers\[53\]\[45\] _10702_ VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__mux2_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _10088_ VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__clkbuf_8
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24881_ _09540_ registers\[53\]\[12\] _10669_ VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__mux2_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26620_ _11622_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23832_ _09644_ registers\[29\]\[62\] _10016_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__mux2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35818_ clknet_leaf_398_CLK _03932_ VGND VGND VPWR VPWR registers\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 _00098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26551_ _11585_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__buf_4
Xclkbuf_5_14_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_14_0_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA_418 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23763_ _09575_ registers\[29\]\[29\] _10039_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__mux2_1
XANTENNA_429 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20975_ _07373_ _07664_ _07665_ _07383_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__a22o_1
XFILLER_122_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35749_ clknet_leaf_462_CLK _03863_ VGND VGND VPWR VPWR registers\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25502_ _11031_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22714_ _07296_ _09353_ _09354_ _07302_ VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__a22o_1
X_29270_ _13079_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__clkbuf_1
X_23694_ registers\[61\]\[62\] _09823_ _09942_ VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__mux2_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26482_ _11549_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28221_ _12496_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22645_ registers\[60\]\[56\] registers\[61\]\[56\] registers\[62\]\[56\] registers\[63\]\[56\]
+ _09227_ _09021_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__mux4_1
X_25433_ _10993_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_179_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_179_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_29_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_29_0_CLK sky130_fd_sc_hd__clkbuf_8
X_28152_ _12460_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__clkbuf_1
X_25364_ _10768_ registers\[50\]\[18\] _10948_ VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22576_ _09155_ _09219_ _09220_ _09158_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__a22o_1
XFILLER_194_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27103_ _11907_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21527_ _08197_ _08201_ _08062_ _08063_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__o211a_1
X_24315_ registers\[57\]\[22\] _10351_ _10347_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__mux2_1
X_28083_ _11843_ registers\[31\]\[54\] _12419_ VGND VGND VPWR VPWR _12424_ sky130_fd_sc_hd__mux2_1
X_25295_ _10864_ VGND VGND VPWR VPWR _10920_ sky130_fd_sc_hd__buf_6
XFILLER_142_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27034_ _11871_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__clkbuf_1
X_24246_ net283 VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21458_ registers\[60\]\[22\] registers\[61\]\[22\] registers\[62\]\[22\] registers\[63\]\[22\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__mux4_1
XFILLER_182_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20409_ registers\[8\]\[58\] registers\[9\]\[58\] registers\[10\]\[58\] registers\[11\]\[58\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__mux4_1
X_24177_ _10268_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_1
X_21389_ registers\[0\]\[20\] registers\[1\]\[20\] registers\[2\]\[20\] registers\[3\]\[20\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_351_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_351_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23128_ registers\[39\]\[13\] _09685_ _09679_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__mux2_1
XTAP_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28985_ _12898_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__clkbuf_1
XTAP_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23059_ net54 VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_103_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_103_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27936_ _12346_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__clkbuf_1
XTAP_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput98 net98 VGND VGND VPWR VPWR D1[17] sky130_fd_sc_hd__buf_2
XTAP_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27867_ _12310_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__clkbuf_1
XTAP_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _04333_ _04401_ _04402_ _04338_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__a22o_1
X_29606_ _13256_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26818_ _11726_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__clkbuf_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27798_ registers\[33\]\[47\] _10403_ _12266_ VGND VGND VPWR VPWR _12274_ sky130_fd_sc_hd__mux2_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29537_ registers\[20\]\[8\] _12951_ _13211_ VGND VGND VPWR VPWR _13220_ sky130_fd_sc_hd__mux2_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ registers\[40\]\[42\] registers\[41\]\[42\] registers\[42\]\[42\] registers\[43\]\[42\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__mux4_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26749_ _11690_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_1
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_930 _09869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ registers\[56\]\[12\] registers\[57\]\[12\] registers\[58\]\[12\] registers\[59\]\[12\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _15004_ sky130_fd_sc_hd__mux4_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_941 _10319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29468_ _13183_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_952 _10439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17482_ _15949_ _15954_ _15955_ VGND VGND VPWR VPWR _15956_ sky130_fd_sc_hd__o21ba_1
XANTENNA_963 _10852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_974 _11158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19221_ registers\[48\]\[24\] registers\[49\]\[24\] registers\[50\]\[24\] registers\[51\]\[24\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__mux4_1
X_28419_ _11774_ registers\[28\]\[21\] _12599_ VGND VGND VPWR VPWR _12601_ sky130_fd_sc_hd__mux2_1
X_16433_ registers\[8\]\[10\] registers\[9\]\[10\] registers\[10\]\[10\] registers\[11\]\[10\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14937_ sky130_fd_sc_hd__mux4_1
XANTENNA_985 _11476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_996 _11795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29399_ _13147_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31430_ _09676_ registers\[6\]\[9\] _14206_ VGND VGND VPWR VPWR _14216_ sky130_fd_sc_hd__mux2_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19152_ _05065_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__buf_4
X_16364_ registers\[8\]\[8\] registers\[9\]\[8\] registers\[10\]\[8\] registers\[11\]\[8\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14870_ sky130_fd_sc_hd__mux4_1
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18103_ registers\[48\]\[58\] registers\[49\]\[58\] registers\[50\]\[58\] registers\[51\]\[58\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__mux4_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19083_ _05102_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__clkbuf_4
X_31361_ registers\[7\]\[40\] net35 _14179_ VGND VGND VPWR VPWR _14180_ sky130_fd_sc_hd__mux2_1
X_16295_ registers\[4\]\[6\] registers\[5\]\[6\] registers\[6\]\[6\] registers\[7\]\[6\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14803_ sky130_fd_sc_hd__mux4_1
XFILLER_240_1290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33100_ clknet_leaf_168_CLK _01214_ VGND VGND VPWR VPWR registers\[51\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30312_ _13627_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__clkbuf_1
X_18034_ _04805_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_2
X_34080_ clknet_leaf_17_CLK _02194_ VGND VGND VPWR VPWR registers\[35\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31292_ _14143_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33031_ clknet_leaf_267_CLK _01145_ VGND VGND VPWR VPWR registers\[52\]\[57\] sky130_fd_sc_hd__dfxtp_2
X_30243_ _13591_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_342_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_342_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30174_ registers\[16\]\[54\] _13048_ _13550_ VGND VGND VPWR VPWR _13555_ sky130_fd_sc_hd__mux2_1
XFILLER_207_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19985_ registers\[32\]\[46\] registers\[33\]\[46\] registers\[34\]\[46\] registers\[35\]\[46\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux4_1
XFILLER_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18936_ _05095_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__clkbuf_8
XFILLER_171_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34982_ clknet_leaf_455_CLK _03096_ VGND VGND VPWR VPWR registers\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1340 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1351 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1362 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33933_ clknet_leaf_168_CLK _02047_ VGND VGND VPWR VPWR registers\[38\]\[63\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1373 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18867_ registers\[56\]\[14\] registers\[57\]\[14\] registers\[58\]\[14\] registers\[59\]\[14\]
+ _05615_ _05405_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__mux4_1
XANTENNA_1384 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1395 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17818_ registers\[16\]\[49\] registers\[17\]\[49\] registers\[18\]\[49\] registers\[19\]\[49\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__mux4_1
X_33864_ clknet_leaf_218_CLK _01978_ VGND VGND VPWR VPWR registers\[3\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18798_ registers\[36\]\[12\] registers\[37\]\[12\] registers\[38\]\[12\] registers\[39\]\[12\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__mux4_1
XFILLER_36_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35603_ clknet_leaf_79_CLK _03717_ VGND VGND VPWR VPWR registers\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_32815_ clknet_leaf_368_CLK _00929_ VGND VGND VPWR VPWR registers\[55\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_17749_ registers\[20\]\[47\] registers\[21\]\[47\] registers\[22\]\[47\] registers\[23\]\[47\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33795_ clknet_leaf_249_CLK _01909_ VGND VGND VPWR VPWR registers\[40\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35534_ clknet_leaf_136_CLK _03648_ VGND VGND VPWR VPWR registers\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_20760_ registers\[4\]\[2\] registers\[5\]\[2\] registers\[6\]\[2\] registers\[7\]\[2\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__mux4_1
XFILLER_63_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32746_ clknet_leaf_420_CLK _00860_ VGND VGND VPWR VPWR registers\[56\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19419_ _06152_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__clkbuf_1
X_35465_ clknet_leaf_159_CLK _03579_ VGND VGND VPWR VPWR registers\[14\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20691_ registers\[28\]\[0\] registers\[29\]\[0\] registers\[30\]\[0\] registers\[31\]\[0\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__mux4_1
X_32677_ clknet_leaf_439_CLK _00791_ VGND VGND VPWR VPWR registers\[57\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22430_ _07333_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__clkbuf_4
X_34416_ clknet_leaf_387_CLK _02530_ VGND VGND VPWR VPWR registers\[30\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_31628_ registers\[63\]\[39\] net33 _14310_ VGND VGND VPWR VPWR _14320_ sky130_fd_sc_hd__mux2_1
X_35396_ clknet_leaf_231_CLK _03510_ VGND VGND VPWR VPWR registers\[15\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22361_ _07274_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__buf_2
XFILLER_17_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34347_ clknet_leaf_401_CLK _02461_ VGND VGND VPWR VPWR registers\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31559_ registers\[63\]\[6\] net61 _14277_ VGND VGND VPWR VPWR _14284_ sky130_fd_sc_hd__mux2_1
X_24100_ _09640_ registers\[5\]\[60\] _10160_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__mux2_1
XFILLER_176_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21312_ registers\[60\]\[18\] registers\[61\]\[18\] registers\[62\]\[18\] registers\[63\]\[18\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__mux4_1
X_25080_ _10790_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
X_22292_ registers\[48\]\[46\] registers\[49\]\[46\] registers\[50\]\[46\] registers\[51\]\[46\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__mux4_1
X_34278_ clknet_leaf_432_CLK _02392_ VGND VGND VPWR VPWR registers\[32\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36017_ clknet_leaf_369_CLK _04131_ VGND VGND VPWR VPWR registers\[63\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_24031_ _09571_ registers\[5\]\[27\] _10183_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__mux2_1
X_33229_ clknet_leaf_144_CLK _01343_ VGND VGND VPWR VPWR registers\[4\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_21243_ registers\[0\]\[16\] registers\[1\]\[16\] registers\[2\]\[16\] registers\[3\]\[16\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_333_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_333_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21174_ _07854_ _07858_ _07719_ _07720_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__o211a_1
XFILLER_171_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20125_ _06838_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
X_28770_ _11855_ registers\[26\]\[60\] _12718_ VGND VGND VPWR VPWR _12785_ sky130_fd_sc_hd__mux2_1
X_25982_ _11286_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27721_ registers\[33\]\[10\] _10325_ _12233_ VGND VGND VPWR VPWR _12234_ sky130_fd_sc_hd__mux2_1
X_20056_ _06569_ _06769_ _06770_ _06574_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__a22o_1
X_24933_ _09592_ registers\[53\]\[37\] _10691_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__mux2_1
XFILLER_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27652_ _12197_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__clkbuf_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24864_ _09523_ registers\[53\]\[4\] _10658_ VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__mux2_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26603_ _11613_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ _10076_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_204 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27583_ registers\[34\]\[9\] _10323_ _12151_ VGND VGND VPWR VPWR _12161_ sky130_fd_sc_hd__mux2_1
XFILLER_26_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24795_ _10626_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_215 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_237 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29322_ _09762_ registers\[22\]\[34\] _13102_ VGND VGND VPWR VPWR _13107_ sky130_fd_sc_hd__mux2_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ _11576_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_248 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20958_ _07328_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_259 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23746_ _10040_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29253_ _09660_ registers\[22\]\[1\] _13069_ VGND VGND VPWR VPWR _13071_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26465_ _11540_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__clkbuf_1
X_23677_ _10002_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
X_20889_ registers\[8\]\[6\] registers\[9\]\[6\] registers\[10\]\[6\] registers\[11\]\[6\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__mux4_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28204_ _12487_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25416_ _10984_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__clkbuf_1
X_22628_ _09104_ _09270_ _09271_ _09107_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__a22o_1
X_29184_ _13024_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__clkbuf_1
X_26396_ _10846_ registers\[43\]\[55\] _11498_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__mux2_1
XFILLER_195_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28135_ _12451_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__clkbuf_1
X_22559_ registers\[4\]\[53\] registers\[5\]\[53\] registers\[6\]\[53\] registers\[7\]\[53\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__mux4_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25347_ _10936_ VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__buf_4
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28066_ _11826_ registers\[31\]\[46\] _12408_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__mux2_1
X_16080_ _14531_ VGND VGND VPWR VPWR _14594_ sky130_fd_sc_hd__buf_12
XFILLER_10_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25278_ _10911_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27017_ net60 VGND VGND VPWR VPWR _11861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24229_ _10295_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_324_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_324_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19770_ _06490_ _06493_ _06194_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o21ba_1
X_28968_ _12889_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__clkbuf_1
X_16982_ registers\[36\]\[26\] registers\[37\]\[26\] registers\[38\]\[26\] registers\[39\]\[26\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15470_ sky130_fd_sc_hd__mux4_1
XFILLER_77_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18721_ _05204_ _05472_ _05473_ _05207_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a22o_1
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27919_ registers\[32\]\[40\] _10388_ _12337_ VGND VGND VPWR VPWR _12338_ sky130_fd_sc_hd__mux2_1
XFILLER_237_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28899_ _11849_ registers\[25\]\[57\] _12845_ VGND VGND VPWR VPWR _12853_ sky130_fd_sc_hd__mux2_1
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _05042_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__buf_4
X_30930_ registers\[10\]\[28\] _12993_ _13944_ VGND VGND VPWR VPWR _13953_ sky130_fd_sc_hd__mux2_1
XFILLER_231_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17603_ _14518_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__buf_6
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30861_ _13916_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__clkbuf_1
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _05095_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__buf_4
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32600_ clknet_leaf_68_CLK _00714_ VGND VGND VPWR VPWR registers\[58\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _15825_ _04318_ _04319_ _15828_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a22o_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33580_ clknet_leaf_330_CLK _01694_ VGND VGND VPWR VPWR registers\[43\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_30792_ _13880_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_760 _07398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32531_ clknet_leaf_78_CLK _00645_ VGND VGND VPWR VPWR registers\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_771 _07890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_782 _08576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17465_ registers\[16\]\[39\] registers\[17\]\[39\] registers\[18\]\[39\] registers\[19\]\[39\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _15940_ sky130_fd_sc_hd__mux4_1
XFILLER_178_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_793 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19204_ registers\[16\]\[23\] registers\[17\]\[23\] registers\[18\]\[23\] registers\[19\]\[23\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__mux4_1
X_16416_ _14648_ _14918_ _14919_ _14653_ VGND VGND VPWR VPWR _14920_ sky130_fd_sc_hd__a22o_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35250_ clknet_leaf_417_CLK _03364_ VGND VGND VPWR VPWR registers\[17\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_32462_ clknet_leaf_178_CLK _00576_ VGND VGND VPWR VPWR registers\[60\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_17396_ registers\[20\]\[37\] registers\[21\]\[37\] registers\[22\]\[37\] registers\[23\]\[37\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15873_ sky130_fd_sc_hd__mux4_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34201_ clknet_leaf_91_CLK _02315_ VGND VGND VPWR VPWR registers\[33\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31413_ _14207_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__clkbuf_1
X_19135_ _05839_ _05875_ _05876_ _05842_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__a22o_1
X_16347_ _14655_ _14851_ _14852_ _14658_ VGND VGND VPWR VPWR _14853_ sky130_fd_sc_hd__a22o_1
X_35181_ clknet_leaf_397_CLK _03295_ VGND VGND VPWR VPWR registers\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_32393_ clknet_leaf_161_CLK _00507_ VGND VGND VPWR VPWR registers\[61\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34132_ clknet_leaf_121_CLK _02246_ VGND VGND VPWR VPWR registers\[34\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31344_ registers\[7\]\[32\] net26 _14168_ VGND VGND VPWR VPWR _14171_ sky130_fd_sc_hd__mux2_1
X_19066_ _05809_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
X_16278_ _14782_ _14785_ _14525_ VGND VGND VPWR VPWR _14786_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18017_ _04548_ _04787_ _04788_ _04552_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a22o_1
X_34063_ clknet_leaf_132_CLK _02177_ VGND VGND VPWR VPWR registers\[35\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31275_ _09656_ _11008_ VGND VGND VPWR VPWR _14134_ sky130_fd_sc_hd__nor2_8
XFILLER_195_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_315_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_315_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_160_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33014_ clknet_leaf_327_CLK _01128_ VGND VGND VPWR VPWR registers\[52\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30226_ _13582_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30157_ registers\[16\]\[46\] _13031_ _13539_ VGND VGND VPWR VPWR _13546_ sky130_fd_sc_hd__mux2_1
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19968_ registers\[8\]\[45\] registers\[9\]\[45\] registers\[10\]\[45\] registers\[11\]\[45\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__mux4_1
XFILLER_101_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18919_ registers\[28\]\[15\] registers\[29\]\[15\] registers\[30\]\[15\] registers\[31\]\[15\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__mux4_1
XFILLER_45_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34965_ clknet_leaf_97_CLK _03079_ VGND VGND VPWR VPWR registers\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1170 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30088_ registers\[16\]\[13\] _12962_ _13506_ VGND VGND VPWR VPWR _13510_ sky130_fd_sc_hd__mux2_1
X_19899_ _06615_ _06618_ _06512_ _06513_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__o211a_1
XFILLER_228_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1181 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1192 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33916_ clknet_leaf_282_CLK _02030_ VGND VGND VPWR VPWR registers\[38\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_21930_ _08593_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__buf_6
XFILLER_83_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34896_ clknet_leaf_115_CLK _03010_ VGND VGND VPWR VPWR registers\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21861_ _08423_ _08525_ _08526_ _08428_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__a22o_1
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33847_ clknet_leaf_316_CLK _01961_ VGND VGND VPWR VPWR registers\[3\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20812_ _07503_ _07506_ _07310_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__o21ba_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ registers\[61\]\[17\] _09693_ _09954_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__mux2_1
XFILLER_242_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24580_ net86 _09649_ net88 VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__and3b_1
XFILLER_110_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21792_ _08456_ _08459_ _08430_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__o21ba_1
X_33778_ clknet_leaf_361_CLK _01892_ VGND VGND VPWR VPWR registers\[40\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23531_ _09924_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
X_35517_ clknet_leaf_297_CLK _03631_ VGND VGND VPWR VPWR registers\[13\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_20743_ _07295_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__buf_6
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32729_ clknet_leaf_68_CLK _00843_ VGND VGND VPWR VPWR registers\[56\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26250_ _11371_ VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23462_ _09888_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20674_ _07372_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__clkbuf_4
X_35448_ clknet_leaf_320_CLK _03562_ VGND VGND VPWR VPWR registers\[14\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22413_ registers\[12\]\[49\] registers\[13\]\[49\] registers\[14\]\[49\] registers\[15\]\[49\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__mux4_1
X_25201_ _10741_ registers\[51\]\[5\] _10865_ VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23393_ _09850_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26181_ _10766_ registers\[44\]\[17\] _11383_ VGND VGND VPWR VPWR _11391_ sky130_fd_sc_hd__mux2_1
X_35379_ clknet_leaf_353_CLK _03493_ VGND VGND VPWR VPWR registers\[15\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22344_ _08992_ _08995_ _08759_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__o21ba_1
X_25132_ _10825_ registers\[52\]\[45\] _10815_ VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29940_ registers\[17\]\[7\] _12949_ _13424_ VGND VGND VPWR VPWR _13432_ sky130_fd_sc_hd__mux2_1
X_25063_ net16 VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_306_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_306_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22275_ registers\[24\]\[45\] registers\[25\]\[45\] registers\[26\]\[45\] registers\[27\]\[45\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__mux4_1
XFILLER_105_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24014_ _09554_ registers\[5\]\[19\] _10172_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__mux2_1
X_21226_ registers\[32\]\[16\] registers\[33\]\[16\] registers\[34\]\[16\] registers\[35\]\[16\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__mux4_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29871_ _13395_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28822_ _11771_ registers\[25\]\[20\] _12812_ VGND VGND VPWR VPWR _12813_ sky130_fd_sc_hd__mux2_1
X_21157_ _07819_ _07826_ _07835_ _07842_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__or4_2
XFILLER_137_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20108_ _06784_ _06820_ _06821_ _06788_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__a22o_1
XFILLER_28_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28753_ _12776_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21088_ _07775_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
X_25965_ _11277_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27704_ registers\[33\]\[2\] _10309_ _12222_ VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__mux2_1
X_20039_ registers\[0\]\[47\] registers\[1\]\[47\] registers\[2\]\[47\] registers\[3\]\[47\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__mux4_1
X_24916_ _09575_ registers\[53\]\[29\] _10680_ VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__mux2_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28684_ _11769_ registers\[26\]\[19\] _12730_ VGND VGND VPWR VPWR _12740_ sky130_fd_sc_hd__mux2_1
XFILLER_218_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25896_ _11229_ VGND VGND VPWR VPWR _11241_ sky130_fd_sc_hd__buf_4
XFILLER_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27635_ _12188_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__clkbuf_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24847_ _10653_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27566_ _12152_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__clkbuf_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _10617_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29305_ _09744_ registers\[22\]\[26\] _13091_ VGND VGND VPWR VPWR _13098_ sky130_fd_sc_hd__mux2_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26517_ _11567_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _10031_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27497_ _11799_ registers\[35\]\[33\] _12111_ VGND VGND VPWR VPWR _12115_ sky130_fd_sc_hd__mux2_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29236_ _13059_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17250_ _14518_ VGND VGND VPWR VPWR _15731_ sky130_fd_sc_hd__buf_6
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26448_ _11531_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16201_ registers\[20\]\[3\] registers\[21\]\[3\] registers\[22\]\[3\] registers\[23\]\[3\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14712_ sky130_fd_sc_hd__mux4_1
XFILLER_122_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17181_ _15482_ _15662_ _15663_ _15485_ VGND VGND VPWR VPWR _15664_ sky130_fd_sc_hd__a22o_1
X_29167_ registers\[23\]\[37\] _13012_ _12998_ VGND VGND VPWR VPWR _13013_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26379_ _10829_ registers\[43\]\[47\] _11487_ VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__mux2_1
XFILLER_35_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16132_ _14601_ _14643_ _14644_ _14611_ VGND VGND VPWR VPWR _14645_ sky130_fd_sc_hd__a22o_1
X_28118_ _12442_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29098_ net7 VGND VGND VPWR VPWR _12966_ sky130_fd_sc_hd__buf_4
X_16063_ _14576_ VGND VGND VPWR VPWR _14577_ sky130_fd_sc_hd__buf_6
XFILLER_170_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28049_ _11809_ registers\[31\]\[38\] _12397_ VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__mux2_1
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31060_ _14021_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30011_ _13469_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19822_ registers\[36\]\[41\] registers\[37\]\[41\] registers\[38\]\[41\] registers\[39\]\[41\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__mux4_1
XFILLER_97_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16965_ registers\[12\]\[25\] registers\[13\]\[25\] registers\[14\]\[25\] registers\[15\]\[25\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15454_ sky130_fd_sc_hd__mux4_1
X_19753_ registers\[60\]\[39\] registers\[61\]\[39\] registers\[62\]\[39\] registers\[63\]\[39\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__mux4_1
XFILLER_46_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18704_ _05454_ _05457_ _05134_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__o21ba_1
XFILLER_42_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34750_ clknet_leaf_179_CLK _02864_ VGND VGND VPWR VPWR registers\[25\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31962_ clknet_leaf_4_CLK _00131_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
X_19684_ _06406_ _06409_ _06169_ _06170_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__o211a_1
XFILLER_231_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16896_ _15139_ _15385_ _15386_ _15142_ VGND VGND VPWR VPWR _15387_ sky130_fd_sc_hd__a22o_1
XFILLER_225_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18635_ _05137_ _05389_ _05390_ _05147_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__a22o_1
X_33701_ clknet_leaf_57_CLK _01815_ VGND VGND VPWR VPWR registers\[41\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_30913_ _13921_ VGND VGND VPWR VPWR _13944_ sky130_fd_sc_hd__buf_4
XFILLER_65_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34681_ clknet_leaf_428_CLK _02795_ VGND VGND VPWR VPWR registers\[26\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31893_ _14459_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33632_ clknet_leaf_33_CLK _01746_ VGND VGND VPWR VPWR registers\[42\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_30844_ _09800_ registers\[11\]\[51\] _13906_ VGND VGND VPWR VPWR _13908_ sky130_fd_sc_hd__mux2_1
X_18566_ registers\[28\]\[5\] registers\[29\]\[5\] registers\[30\]\[5\] registers\[31\]\[5\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__mux4_1
XFILLER_18_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17517_ _04303_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__clkbuf_4
X_33563_ clknet_leaf_26_CLK _01677_ VGND VGND VPWR VPWR registers\[43\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18497_ registers\[24\]\[3\] registers\[25\]\[3\] registers\[26\]\[3\] registers\[27\]\[3\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__mux4_1
X_30775_ _13871_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_590 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32514_ clknet_leaf_201_CLK _00628_ VGND VGND VPWR VPWR registers\[60\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_35302_ clknet_leaf_449_CLK _03416_ VGND VGND VPWR VPWR registers\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17448_ _15684_ _15921_ _15922_ _15687_ VGND VGND VPWR VPWR _15923_ sky130_fd_sc_hd__a22o_1
X_33494_ clknet_leaf_126_CLK _01608_ VGND VGND VPWR VPWR registers\[44\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32445_ clknet_leaf_187_CLK _00559_ VGND VGND VPWR VPWR registers\[29\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_35233_ clknet_leaf_479_CLK _03347_ VGND VGND VPWR VPWR registers\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17379_ registers\[48\]\[37\] registers\[49\]\[37\] registers\[50\]\[37\] registers\[51\]\[37\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15856_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_92_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_92_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19118_ _05856_ _05859_ _05818_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__o21ba_1
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35164_ clknet_leaf_5_CLK _03278_ VGND VGND VPWR VPWR registers\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_20390_ registers\[20\]\[57\] registers\[21\]\[57\] registers\[22\]\[57\] registers\[23\]\[57\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__mux4_1
X_32376_ clknet_leaf_331_CLK _00490_ VGND VGND VPWR VPWR registers\[61\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34115_ clknet_leaf_247_CLK _02229_ VGND VGND VPWR VPWR registers\[35\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31327_ registers\[7\]\[24\] net17 _14157_ VGND VGND VPWR VPWR _14162_ sky130_fd_sc_hd__mux2_1
X_19049_ _05755_ _05791_ _05792_ _05759_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__a22o_1
X_35095_ clknet_leaf_81_CLK _03209_ VGND VGND VPWR VPWR registers\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xoutput200 net200 VGND VGND VPWR VPWR D2[51] sky130_fd_sc_hd__buf_2
XFILLER_133_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput211 net211 VGND VGND VPWR VPWR D2[61] sky130_fd_sc_hd__buf_2
Xoutput222 net222 VGND VGND VPWR VPWR D3[13] sky130_fd_sc_hd__buf_2
X_34046_ clknet_leaf_269_CLK _02160_ VGND VGND VPWR VPWR registers\[36\]\[48\] sky130_fd_sc_hd__dfxtp_1
Xoutput233 net233 VGND VGND VPWR VPWR D3[23] sky130_fd_sc_hd__buf_2
X_22060_ registers\[12\]\[39\] registers\[13\]\[39\] registers\[14\]\[39\] registers\[15\]\[39\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__mux4_1
X_31258_ _14125_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__clkbuf_1
Xoutput244 net244 VGND VGND VPWR VPWR D3[33] sky130_fd_sc_hd__buf_2
Xoutput255 net255 VGND VGND VPWR VPWR D3[43] sky130_fd_sc_hd__buf_2
X_21011_ _07697_ _07700_ _07399_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__o21ba_1
Xoutput266 net266 VGND VGND VPWR VPWR D3[53] sky130_fd_sc_hd__buf_2
XFILLER_82_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30209_ _13573_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput277 net277 VGND VGND VPWR VPWR D3[63] sky130_fd_sc_hd__buf_2
XFILLER_47_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31189_ _14089_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35997_ clknet_leaf_55_CLK _04111_ VGND VGND VPWR VPWR registers\[63\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_25750_ _11164_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
X_34948_ clknet_leaf_202_CLK _03062_ VGND VGND VPWR VPWR registers\[22\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22962_ _09570_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_845 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24701_ _09632_ registers\[55\]\[56\] _10569_ VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__mux2_1
X_21913_ _07287_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__buf_6
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25681_ registers\[48\]\[37\] _10382_ _11119_ VGND VGND VPWR VPWR _11127_ sky130_fd_sc_hd__mux2_1
XFILLER_55_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22893_ _09523_ registers\[62\]\[4\] _09515_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__mux2_1
X_34879_ clknet_leaf_307_CLK _02993_ VGND VGND VPWR VPWR registers\[23\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27420_ registers\[36\]\[61\] _10432_ _12006_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__mux2_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24632_ _09563_ registers\[55\]\[23\] _10536_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__mux2_1
XFILLER_71_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21844_ registers\[52\]\[33\] registers\[53\]\[33\] registers\[54\]\[33\] registers\[55\]\[33\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__mux4_1
XFILLER_215_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27351_ registers\[36\]\[28\] _10363_ _12029_ VGND VGND VPWR VPWR _12038_ sky130_fd_sc_hd__mux2_1
X_24563_ _09632_ registers\[56\]\[56\] _10495_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__mux2_1
XFILLER_196_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21775_ registers\[60\]\[31\] registers\[61\]\[31\] registers\[62\]\[31\] registers\[63\]\[31\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__mux4_1
XFILLER_93_1255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26302_ _10751_ registers\[43\]\[10\] _11454_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__mux2_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20726_ _07420_ _07423_ _07370_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__o21ba_1
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23514_ _09601_ registers\[19\]\[41\] _09914_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__mux2_1
X_27282_ _12001_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24494_ _09563_ registers\[56\]\[23\] _10462_ VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29021_ _12917_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__clkbuf_1
X_26233_ _11418_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
X_20657_ _07277_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__buf_12
X_23445_ _09879_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_83_CLK sky130_fd_sc_hd__clkbuf_16
X_26164_ _10749_ registers\[44\]\[9\] _11372_ VGND VGND VPWR VPWR _11382_ sky130_fd_sc_hd__mux2_1
XFILLER_176_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23376_ registers\[39\]\[41\] _09778_ _09840_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__mux2_1
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20588_ _07277_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__buf_12
XFILLER_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25115_ net35 VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__buf_2
X_22327_ _07358_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__buf_4
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26095_ _10814_ registers\[45\]\[40\] _11345_ VGND VGND VPWR VPWR _11346_ sky130_fd_sc_hd__mux2_1
X_29923_ _13422_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__clkbuf_1
X_22258_ _08908_ _08911_ _08740_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__o21ba_1
X_25046_ _10767_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21209_ registers\[8\]\[15\] registers\[9\]\[15\] registers\[10\]\[15\] registers\[11\]\[15\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__mux4_1
X_29854_ registers\[18\]\[30\] _12997_ _13386_ VGND VGND VPWR VPWR _13387_ sky130_fd_sc_hd__mux2_1
X_22189_ registers\[44\]\[43\] registers\[45\]\[43\] registers\[46\]\[43\] registers\[47\]\[43\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__mux4_1
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28805_ _11755_ registers\[25\]\[12\] _12801_ VGND VGND VPWR VPWR _12804_ sky130_fd_sc_hd__mux2_1
X_29785_ registers\[1\]\[62\] _13064_ _13281_ VGND VGND VPWR VPWR _13350_ sky130_fd_sc_hd__mux2_1
X_26997_ _11847_ registers\[3\]\[56\] _11835_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__mux2_1
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28736_ _12767_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16750_ _15241_ _15244_ _14934_ _14935_ VGND VGND VPWR VPWR _15245_ sky130_fd_sc_hd__o211a_1
XFILLER_47_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25948_ _11268_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16681_ _15139_ _15176_ _15177_ _15142_ VGND VGND VPWR VPWR _15178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28667_ _12731_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__clkbuf_1
X_25879_ _11232_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
X_18420_ registers\[8\]\[1\] registers\[9\]\[1\] registers\[10\]\[1\] registers\[11\]\[1\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__mux4_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27618_ _12179_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28598_ _11818_ registers\[27\]\[42\] _12692_ VGND VGND VPWR VPWR _12695_ sky130_fd_sc_hd__mux2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__clkbuf_4
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27549_ _11851_ registers\[35\]\[58\] _12133_ VGND VGND VPWR VPWR _12142_ sky130_fd_sc_hd__mux2_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ registers\[44\]\[35\] registers\[45\]\[35\] registers\[46\]\[35\] registers\[47\]\[35\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15781_ sky130_fd_sc_hd__mux4_1
XFILLER_230_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__buf_12
X_30560_ _13758_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29219_ net50 VGND VGND VPWR VPWR _13048_ sky130_fd_sc_hd__clkbuf_4
X_17233_ registers\[40\]\[33\] registers\[41\]\[33\] registers\[42\]\[33\] registers\[43\]\[33\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15714_ sky130_fd_sc_hd__mux4_1
XFILLER_202_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30491_ _13722_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_74_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_74_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32230_ clknet_leaf_157_CLK _00344_ VGND VGND VPWR VPWR registers\[9\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17164_ _15647_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16115_ _14528_ _14626_ _14627_ _14537_ VGND VGND VPWR VPWR _14628_ sky130_fd_sc_hd__a22o_1
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32161_ clknet_leaf_40_CLK _00275_ VGND VGND VPWR VPWR registers\[39\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17095_ _15341_ _15578_ _15579_ _15344_ VGND VGND VPWR VPWR _15580_ sky130_fd_sc_hd__a22o_1
XFILLER_182_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31112_ registers\[0\]\[50\] _13039_ _14048_ VGND VGND VPWR VPWR _14049_ sky130_fd_sc_hd__mux2_1
X_16046_ _14504_ VGND VGND VPWR VPWR _14560_ sky130_fd_sc_hd__buf_6
X_32092_ clknet_leaf_489_CLK _00005_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35920_ clknet_leaf_108_CLK _04034_ VGND VGND VPWR VPWR registers\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_31043_ _14012_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19805_ _05116_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35851_ clknet_leaf_151_CLK _03965_ VGND VGND VPWR VPWR registers\[8\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17997_ registers\[16\]\[54\] registers\[17\]\[54\] registers\[18\]\[54\] registers\[19\]\[54\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux4_1
XFILLER_97_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34802_ clknet_leaf_384_CLK _02916_ VGND VGND VPWR VPWR registers\[24\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19736_ registers\[20\]\[38\] registers\[21\]\[38\] registers\[22\]\[38\] registers\[23\]\[38\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__mux4_1
X_16948_ _15334_ _15435_ _15436_ _15339_ VGND VGND VPWR VPWR _15437_ sky130_fd_sc_hd__a22o_1
X_35782_ clknet_leaf_217_CLK _03896_ VGND VGND VPWR VPWR registers\[0\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32994_ clknet_leaf_443_CLK _01108_ VGND VGND VPWR VPWR registers\[52\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34733_ clknet_leaf_410_CLK _02847_ VGND VGND VPWR VPWR registers\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31945_ _14486_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__clkbuf_1
X_19667_ _06364_ _06373_ _06384_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or4_2
X_16879_ _15370_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18618_ _05368_ _05373_ _05074_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19598_ _06326_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__buf_2
X_34664_ clknet_leaf_453_CLK _02778_ VGND VGND VPWR VPWR registers\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31876_ _14450_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33615_ clknet_leaf_131_CLK _01729_ VGND VGND VPWR VPWR registers\[42\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_30827_ _09782_ registers\[11\]\[43\] _13895_ VGND VGND VPWR VPWR _13899_ sky130_fd_sc_hd__mux2_1
X_18549_ _05077_ _05305_ _05306_ _05086_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__a22o_1
XFILLER_212_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34595_ clknet_leaf_445_CLK _02709_ VGND VGND VPWR VPWR registers\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21560_ _07287_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__buf_4
X_33546_ clknet_leaf_162_CLK _01660_ VGND VGND VPWR VPWR registers\[44\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30758_ _09678_ registers\[11\]\[10\] _13862_ VGND VGND VPWR VPWR _13863_ sky130_fd_sc_hd__mux2_1
X_20511_ _05119_ _07211_ _07212_ _05131_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__a22o_1
XFILLER_127_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33477_ clknet_leaf_255_CLK _01591_ VGND VGND VPWR VPWR registers\[45\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_21491_ registers\[52\]\[23\] registers\[53\]\[23\] registers\[54\]\[23\] registers\[55\]\[23\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_65_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_65_CLK sky130_fd_sc_hd__clkbuf_16
X_30689_ _13826_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23230_ _09748_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
X_20442_ registers\[12\]\[59\] registers\[13\]\[59\] registers\[14\]\[59\] registers\[15\]\[59\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__mux4_1
X_35216_ clknet_leaf_114_CLK _03330_ VGND VGND VPWR VPWR registers\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_32428_ clknet_leaf_396_CLK _00542_ VGND VGND VPWR VPWR registers\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36196_ clknet_leaf_92_CLK _00078_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23161_ registers\[9\]\[0\] _09648_ _09709_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__mux2_1
X_35147_ clknet_leaf_151_CLK _03261_ VGND VGND VPWR VPWR registers\[1\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_20373_ registers\[48\]\[57\] registers\[49\]\[57\] registers\[50\]\[57\] registers\[51\]\[57\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__mux4_1
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32359_ clknet_leaf_436_CLK _00473_ VGND VGND VPWR VPWR registers\[61\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22112_ _07366_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__clkbuf_4
XTAP_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23092_ _09661_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
X_35078_ clknet_leaf_208_CLK _03192_ VGND VGND VPWR VPWR registers\[20\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22043_ _07305_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__buf_4
X_26920_ _11795_ registers\[3\]\[31\] _11793_ VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__mux2_1
X_34029_ clknet_leaf_327_CLK _02143_ VGND VGND VPWR VPWR registers\[36\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26851_ _11748_ registers\[3\]\[9\] _11730_ VGND VGND VPWR VPWR _11749_ sky130_fd_sc_hd__mux2_1
XFILLER_141_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25802_ _11191_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
X_29570_ _13237_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26782_ registers\[40\]\[45\] _10399_ _11702_ VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__mux2_1
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23994_ _10171_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28521_ _12654_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__clkbuf_1
X_25733_ registers\[48\]\[62\] _10434_ _11085_ VGND VGND VPWR VPWR _11154_ sky130_fd_sc_hd__mux2_1
X_22945_ net14 VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__buf_2
XFILLER_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28452_ _11807_ registers\[28\]\[37\] _12610_ VGND VGND VPWR VPWR _12618_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25664_ registers\[48\]\[29\] _10365_ _11108_ VGND VGND VPWR VPWR _11118_ sky130_fd_sc_hd__mux2_1
X_22876_ net85 net84 VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__nand2_8
XFILLER_147_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27403_ _12065_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24615_ _09546_ registers\[55\]\[15\] _10525_ VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__mux2_1
XFILLER_227_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28383_ _11738_ registers\[28\]\[4\] _12577_ VGND VGND VPWR VPWR _12582_ sky130_fd_sc_hd__mux2_1
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21827_ registers\[28\]\[32\] registers\[29\]\[32\] registers\[30\]\[32\] registers\[31\]\[32\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__mux4_1
X_25595_ registers\[4\]\[62\] _10434_ _11011_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__mux2_1
XFILLER_12_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27334_ _12006_ VGND VGND VPWR VPWR _12029_ sky130_fd_sc_hd__buf_4
XFILLER_223_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24546_ _09615_ registers\[56\]\[48\] _10484_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21758_ registers\[20\]\[30\] registers\[21\]\[30\] registers\[22\]\[30\] registers\[23\]\[30\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__mux4_1
XFILLER_223_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20709_ _07358_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__buf_4
XFILLER_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27265_ _11837_ registers\[37\]\[51\] _11991_ VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__mux2_1
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24477_ _09546_ registers\[56\]\[15\] _10451_ VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__mux2_1
X_21689_ _07303_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_56_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_56_CLK sky130_fd_sc_hd__clkbuf_16
X_29004_ _12908_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__clkbuf_1
X_26216_ _11409_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
X_23428_ _09510_ registers\[19\]\[0\] _09870_ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__mux2_1
XFILLER_149_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27196_ _11956_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26147_ _11373_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23359_ registers\[39\]\[33\] _09760_ _09829_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__mux2_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26078_ _10798_ registers\[45\]\[32\] _11334_ VGND VGND VPWR VPWR _11337_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29906_ registers\[18\]\[55\] _13050_ _13408_ VGND VGND VPWR VPWR _13414_ sky130_fd_sc_hd__mux2_1
X_17920_ _04691_ _04694_ _04619_ _04620_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__o211a_1
X_25029_ net4 VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__clkbuf_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1703 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1714 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1725 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1736 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17851_ registers\[4\]\[50\] registers\[5\]\[50\] registers\[6\]\[50\] registers\[7\]\[50\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__mux4_1
XTAP_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1747 _05067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29837_ registers\[18\]\[22\] _12981_ _13375_ VGND VGND VPWR VPWR _13378_ sky130_fd_sc_hd__mux2_1
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1758 _07338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_45__f_CLK clknet_5_22_0_CLK VGND VGND VPWR VPWR clknet_6_45__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1769 _09666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16802_ registers\[28\]\[20\] registers\[29\]\[20\] registers\[30\]\[20\] registers\[31\]\[20\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15296_ sky130_fd_sc_hd__mux4_1
XTAP_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17782_ registers\[4\]\[48\] registers\[5\]\[48\] registers\[6\]\[48\] registers\[7\]\[48\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__mux4_1
X_29768_ _13341_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19521_ _06248_ _06251_ _06180_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__o21ba_1
X_16733_ _15197_ _15212_ _15221_ _15228_ VGND VGND VPWR VPWR _15229_ sky130_fd_sc_hd__or4_1
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28719_ _12758_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__clkbuf_1
X_29699_ _13305_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19452_ _05146_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__clkbuf_4
X_31730_ registers\[59\]\[23\] net16 _14370_ VGND VGND VPWR VPWR _14374_ sky130_fd_sc_hd__mux2_1
XFILLER_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16664_ registers\[32\]\[17\] registers\[33\]\[17\] registers\[34\]\[17\] registers\[35\]\[17\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15161_ sky130_fd_sc_hd__mux4_1
XFILLER_234_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18403_ _05165_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31661_ _14337_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__clkbuf_1
X_19383_ registers\[20\]\[28\] registers\[21\]\[28\] registers\[22\]\[28\] registers\[23\]\[28\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__mux4_1
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16595_ _14991_ _15092_ _15093_ _14996_ VGND VGND VPWR VPWR _15094_ sky130_fd_sc_hd__a22o_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18334_ _05044_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__buf_12
X_30612_ registers\[12\]\[5\] _12945_ _13780_ VGND VGND VPWR VPWR _13786_ sky130_fd_sc_hd__mux2_1
X_33400_ clknet_leaf_340_CLK _01514_ VGND VGND VPWR VPWR registers\[46\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_34380_ clknet_leaf_140_CLK _02494_ VGND VGND VPWR VPWR registers\[31\]\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31592_ _14301_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33331_ clknet_leaf_346_CLK _01445_ VGND VGND VPWR VPWR registers\[47\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_18265_ _05025_ _05028_ _14584_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__o21ba_1
XFILLER_203_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30543_ _13749_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_47_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17216_ registers\[0\]\[32\] registers\[1\]\[32\] registers\[2\]\[32\] registers\[3\]\[32\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15698_ sky130_fd_sc_hd__mux4_1
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36050_ clknet_leaf_71_CLK _04164_ VGND VGND VPWR VPWR registers\[59\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33262_ clknet_leaf_365_CLK _01376_ VGND VGND VPWR VPWR registers\[48\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_18196_ registers\[52\]\[61\] registers\[53\]\[61\] registers\[54\]\[61\] registers\[55\]\[61\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__mux4_1
X_30474_ _13713_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32213_ clknet_leaf_288_CLK _00327_ VGND VGND VPWR VPWR registers\[9\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35001_ clknet_leaf_308_CLK _03115_ VGND VGND VPWR VPWR registers\[21\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17147_ _14584_ VGND VGND VPWR VPWR _15631_ sky130_fd_sc_hd__clkbuf_4
X_33193_ clknet_leaf_401_CLK _01307_ VGND VGND VPWR VPWR registers\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32144_ clknet_leaf_135_CLK _00258_ VGND VGND VPWR VPWR registers\[39\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_17078_ _15558_ _15563_ _15288_ VGND VGND VPWR VPWR _15564_ sky130_fd_sc_hd__o21ba_1
XFILLER_226_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16029_ _14495_ VGND VGND VPWR VPWR _14543_ sky130_fd_sc_hd__buf_12
X_32075_ clknet_leaf_167_CLK _00253_ VGND VGND VPWR VPWR registers\[62\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35903_ clknet_leaf_295_CLK _04017_ VGND VGND VPWR VPWR registers\[7\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_31026_ _14003_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35834_ clknet_leaf_332_CLK _03948_ VGND VGND VPWR VPWR registers\[8\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_19719_ registers\[52\]\[38\] registers\[53\]\[38\] registers\[54\]\[38\] registers\[55\]\[38\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__mux4_1
X_20991_ registers\[56\]\[9\] registers\[57\]\[9\] registers\[58\]\[9\] registers\[59\]\[9\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__mux4_1
X_35765_ clknet_leaf_354_CLK _03879_ VGND VGND VPWR VPWR registers\[0\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32977_ clknet_leaf_173_CLK _01091_ VGND VGND VPWR VPWR registers\[52\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22730_ _09155_ _09368_ _09369_ _09158_ VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__a22o_1
X_34716_ clknet_leaf_5_CLK _02830_ VGND VGND VPWR VPWR registers\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_31928_ _09804_ registers\[49\]\[53\] _14474_ VGND VGND VPWR VPWR _14478_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35696_ clknet_leaf_376_CLK _03810_ VGND VGND VPWR VPWR registers\[10\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22661_ _09109_ _09302_ _09303_ _09114_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__a22o_1
X_34647_ clknet_leaf_93_CLK _02761_ VGND VGND VPWR VPWR registers\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31859_ _09699_ registers\[49\]\[20\] _14441_ VGND VGND VPWR VPWR _14442_ sky130_fd_sc_hd__mux2_1
X_24400_ net46 VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__buf_4
XFILLER_209_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21612_ _08080_ _08283_ _08284_ _08085_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__a22o_1
XFILLER_55_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25380_ _10965_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__clkbuf_1
X_22592_ _08958_ _09235_ _09236_ _08961_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__a22o_1
X_34578_ clknet_leaf_95_CLK _02692_ VGND VGND VPWR VPWR registers\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24331_ _10362_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33529_ clknet_leaf_339_CLK _01643_ VGND VGND VPWR VPWR registers\[44\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_21543_ _08214_ _08217_ _08087_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__o21ba_1
XFILLER_181_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_38_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_38_CLK sky130_fd_sc_hd__clkbuf_16
X_27050_ _11757_ registers\[38\]\[13\] _11876_ VGND VGND VPWR VPWR _11880_ sky130_fd_sc_hd__mux2_1
X_24262_ registers\[57\]\[5\] _10315_ _10305_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__mux2_1
X_21474_ registers\[28\]\[22\] registers\[29\]\[22\] registers\[30\]\[22\] registers\[31\]\[22\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__mux4_1
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26001_ _10856_ registers\[46\]\[60\] _11229_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__mux2_1
XFILLER_140_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20425_ registers\[40\]\[59\] registers\[41\]\[59\] registers\[42\]\[59\] registers\[43\]\[59\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__mux4_1
X_23213_ registers\[9\]\[22\] _09717_ _09735_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__mux2_1
XFILLER_181_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36179_ clknet_leaf_93_CLK _00119_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dfxtp_1
X_24193_ _10276_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20356_ registers\[24\]\[56\] registers\[25\]\[56\] registers\[26\]\[56\] registers\[27\]\[56\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__mux4_1
X_23144_ _09696_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XTAP_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27952_ registers\[32\]\[56\] _10422_ _12348_ VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__mux2_1
X_23075_ _09646_ registers\[62\]\[63\] _09514_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__mux2_1
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20287_ registers\[8\]\[54\] registers\[9\]\[54\] registers\[10\]\[54\] registers\[11\]\[54\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__mux4_1
XTAP_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26903_ net19 VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__buf_2
XFILLER_66_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22026_ registers\[12\]\[38\] registers\[13\]\[38\] registers\[14\]\[38\] registers\[15\]\[38\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__mux4_1
XTAP_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27883_ registers\[32\]\[23\] _10353_ _12315_ VGND VGND VPWR VPWR _12319_ sky130_fd_sc_hd__mux2_1
XFILLER_212_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26834_ _11737_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29622_ _13264_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29553_ _13228_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__clkbuf_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26765_ registers\[40\]\[37\] _10382_ _11691_ VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__mux2_1
X_23977_ _09517_ registers\[5\]\[1\] _10161_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__mux2_1
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28504_ _11859_ registers\[28\]\[62\] _12576_ VGND VGND VPWR VPWR _12645_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25716_ _11145_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29484_ _09791_ registers\[21\]\[47\] _13184_ VGND VGND VPWR VPWR _13192_ sky130_fd_sc_hd__mux2_1
X_22928_ _09547_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26696_ registers\[40\]\[4\] _10313_ _11658_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__mux2_1
XFILLER_16_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28435_ _11790_ registers\[28\]\[29\] _12599_ VGND VGND VPWR VPWR _12609_ sky130_fd_sc_hd__mux2_1
XFILLER_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25647_ _11109_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
X_22859_ registers\[8\]\[63\] registers\[9\]\[63\] registers\[10\]\[63\] registers\[11\]\[63\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__mux4_1
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28366_ _12572_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__clkbuf_1
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _14854_ _14869_ _14878_ _14885_ VGND VGND VPWR VPWR _14886_ sky130_fd_sc_hd__or4_4
X_25578_ _11071_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27317_ _12020_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24529_ _10439_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__buf_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28297_ _12536_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__clkbuf_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_29_CLK sky130_fd_sc_hd__clkbuf_16
X_18050_ registers\[0\]\[56\] registers\[1\]\[56\] registers\[2\]\[56\] registers\[3\]\[56\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__mux4_1
XFILLER_240_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27248_ _11820_ registers\[37\]\[43\] _11980_ VGND VGND VPWR VPWR _11984_ sky130_fd_sc_hd__mux2_1
XFILLER_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17001_ registers\[4\]\[26\] registers\[5\]\[26\] registers\[6\]\[26\] registers\[7\]\[26\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15489_ sky130_fd_sc_hd__mux4_1
XFILLER_158_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27179_ _11750_ registers\[37\]\[10\] _11947_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30190_ registers\[16\]\[62\] _13064_ _13494_ VGND VGND VPWR VPWR _13563_ sky130_fd_sc_hd__mux2_1
XFILLER_126_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18952_ registers\[24\]\[16\] registers\[25\]\[16\] registers\[26\]\[16\] registers\[27\]\[16\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__mux4_1
XANTENNA_1500 _07333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1511 _07507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1522 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17903_ _14496_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__buf_6
XANTENNA_1533 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1544 _10232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18883_ _05113_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__buf_4
XTAP_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1555 _11513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1566 _11935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32900_ clknet_leaf_199_CLK _01014_ VGND VGND VPWR VPWR registers\[54\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17834_ _14524_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__buf_2
XFILLER_66_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1577 _13708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1588 _14493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33880_ clknet_leaf_31_CLK _01994_ VGND VGND VPWR VPWR registers\[38\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1599 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32831_ clknet_leaf_292_CLK _00945_ VGND VGND VPWR VPWR registers\[55\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_17765_ _14543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19504_ registers\[36\]\[32\] registers\[37\]\[32\] registers\[38\]\[32\] registers\[39\]\[32\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__mux4_1
X_35550_ clknet_leaf_484_CLK _03664_ VGND VGND VPWR VPWR registers\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_16716_ _15205_ _15211_ _14934_ _14935_ VGND VGND VPWR VPWR _15212_ sky130_fd_sc_hd__o211a_1
XFILLER_78_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17696_ _14548_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__clkbuf_4
X_32762_ clknet_leaf_284_CLK _00876_ VGND VGND VPWR VPWR registers\[56\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34501_ clknet_leaf_226_CLK _02615_ VGND VGND VPWR VPWR registers\[2\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19435_ _06098_ _06166_ _06167_ _06102_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__a22o_1
X_16647_ registers\[12\]\[16\] registers\[13\]\[16\] registers\[14\]\[16\] registers\[15\]\[16\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15145_ sky130_fd_sc_hd__mux4_1
X_31713_ registers\[59\]\[15\] net7 _14359_ VGND VGND VPWR VPWR _14365_ sky130_fd_sc_hd__mux2_1
X_35481_ clknet_leaf_43_CLK _03595_ VGND VGND VPWR VPWR registers\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_32693_ clknet_leaf_351_CLK _00807_ VGND VGND VPWR VPWR registers\[57\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34432_ clknet_leaf_199_CLK _02546_ VGND VGND VPWR VPWR registers\[30\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_31644_ _14328_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__clkbuf_1
X_16578_ registers\[12\]\[14\] registers\[13\]\[14\] registers\[14\]\[14\] registers\[15\]\[14\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15078_ sky130_fd_sc_hd__mux4_1
XFILLER_37_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19366_ registers\[52\]\[28\] registers\[53\]\[28\] registers\[54\]\[28\] registers\[55\]\[28\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__mux4_1
XFILLER_210_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18317_ _05044_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__buf_12
X_34363_ clknet_leaf_184_CLK _02477_ VGND VGND VPWR VPWR registers\[31\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_31575_ _14292_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__clkbuf_1
X_19297_ _05116_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36102_ clknet_leaf_261_CLK _04216_ VGND VGND VPWR VPWR registers\[59\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18248_ registers\[44\]\[63\] registers\[45\]\[63\] registers\[46\]\[63\] registers\[47\]\[63\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__mux4_1
XFILLER_148_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33314_ clknet_leaf_58_CLK _01428_ VGND VGND VPWR VPWR registers\[47\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_30526_ _13740_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__clkbuf_1
X_34294_ clknet_leaf_341_CLK _02408_ VGND VGND VPWR VPWR registers\[32\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36033_ clknet_leaf_265_CLK _04147_ VGND VGND VPWR VPWR registers\[63\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30457_ _09819_ registers\[14\]\[60\] _13637_ VGND VGND VPWR VPWR _13704_ sky130_fd_sc_hd__mux2_1
X_18179_ registers\[28\]\[60\] registers\[29\]\[60\] registers\[30\]\[60\] registers\[31\]\[60\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__mux4_1
XFILLER_163_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33245_ clknet_leaf_51_CLK _01359_ VGND VGND VPWR VPWR registers\[48\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20210_ registers\[36\]\[52\] registers\[37\]\[52\] registers\[38\]\[52\] registers\[39\]\[52\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux4_1
XFILLER_128_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33176_ clknet_leaf_474_CLK _01290_ VGND VGND VPWR VPWR registers\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_21190_ _07871_ _07874_ _07744_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__o21ba_1
X_30388_ _09747_ registers\[14\]\[27\] _13660_ VGND VGND VPWR VPWR _13668_ sky130_fd_sc_hd__mux2_1
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20141_ _06784_ _06852_ _06853_ _06788_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__a22o_1
XFILLER_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32127_ clknet_leaf_393_CLK _00043_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20072_ registers\[52\]\[48\] registers\[53\]\[48\] registers\[54\]\[48\] registers\[55\]\[48\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__mux4_1
X_32058_ clknet_leaf_287_CLK _00236_ VGND VGND VPWR VPWR registers\[62\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31009_ registers\[0\]\[1\] _12937_ _13993_ VGND VGND VPWR VPWR _13995_ sky130_fd_sc_hd__mux2_1
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23900_ _10121_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24880_ _10671_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23831_ _10084_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__clkbuf_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35817_ clknet_leaf_399_CLK _03931_ VGND VGND VPWR VPWR registers\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26550_ _11584_ _11157_ VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__nand2_8
XANTENNA_408 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35748_ clknet_leaf_465_CLK _03862_ VGND VGND VPWR VPWR registers\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_23762_ _10048_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ registers\[16\]\[8\] registers\[17\]\[8\] registers\[18\]\[8\] registers\[19\]\[8\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__mux4_1
XANTENNA_419 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25501_ registers\[4\]\[17\] _10340_ _11023_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__mux2_1
XFILLER_96_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22713_ registers\[4\]\[58\] registers\[5\]\[58\] registers\[6\]\[58\] registers\[7\]\[58\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__mux4_1
XFILLER_198_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26481_ _10796_ registers\[42\]\[31\] _11547_ VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23693_ _10010_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
X_35679_ clknet_leaf_488_CLK _03793_ VGND VGND VPWR VPWR registers\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28220_ _11845_ registers\[30\]\[55\] _12490_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25432_ _10835_ registers\[50\]\[50\] _10992_ VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__mux2_1
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22644_ _09012_ _09285_ _09286_ _09018_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__a22o_1
XFILLER_55_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28151_ _11776_ registers\[30\]\[22\] _12457_ VGND VGND VPWR VPWR _12460_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25363_ _10956_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__clkbuf_1
X_22575_ registers\[36\]\[54\] registers\[37\]\[54\] registers\[38\]\[54\] registers\[39\]\[54\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_9__f_CLK clknet_5_4_0_CLK VGND VGND VPWR VPWR clknet_6_9__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27102_ _11809_ registers\[38\]\[38\] _11898_ VGND VGND VPWR VPWR _11907_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24314_ net15 VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__clkbuf_4
X_28082_ _12423_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__clkbuf_1
X_21526_ _07991_ _08199_ _08200_ _07995_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__a22o_1
XFILLER_107_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25294_ _10919_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27033_ _11740_ registers\[38\]\[5\] _11865_ VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24245_ net85 net84 _09940_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__nor3_4
X_21457_ _07983_ _08132_ _08133_ _07989_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__a22o_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20408_ _07109_ _07112_ _06855_ _06856_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__o211a_1
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24176_ _09580_ registers\[58\]\[31\] _10266_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__mux2_1
X_21388_ _07349_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23127_ net5 VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__buf_6
X_20339_ registers\[36\]\[56\] registers\[37\]\[56\] registers\[38\]\[56\] registers\[39\]\[56\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__mux4_1
XTAP_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28984_ registers\[24\]\[33\] _10374_ _12894_ VGND VGND VPWR VPWR _12898_ sky130_fd_sc_hd__mux2_1
XTAP_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23058_ _09635_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27935_ registers\[32\]\[48\] _10405_ _12337_ VGND VGND VPWR VPWR _12346_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 net99 VGND VGND VPWR VPWR D1[18] sky130_fd_sc_hd__buf_2
XTAP_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22009_ _07316_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__buf_4
XTAP_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27866_ registers\[32\]\[15\] _10336_ _12304_ VGND VGND VPWR VPWR _12310_ sky130_fd_sc_hd__mux2_1
XFILLER_248_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29605_ registers\[20\]\[40\] _13018_ _13255_ VGND VGND VPWR VPWR _13256_ sky130_fd_sc_hd__mux2_1
X_26817_ registers\[40\]\[62\] _10434_ _11657_ VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__mux2_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27797_ _12273_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__clkbuf_1
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17550_ _14496_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__clkbuf_4
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29536_ _13219_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__clkbuf_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26748_ registers\[40\]\[29\] _10365_ _11680_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__mux2_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16501_ _14997_ _15002_ _14926_ VGND VGND VPWR VPWR _15003_ sky130_fd_sc_hd__o21ba_1
XANTENNA_920 _09778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_931 _09942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29467_ _09773_ registers\[21\]\[39\] _13173_ VGND VGND VPWR VPWR _13183_ sky130_fd_sc_hd__mux2_1
XANTENNA_942 _10328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17481_ _14524_ VGND VGND VPWR VPWR _15955_ sky130_fd_sc_hd__buf_2
X_26679_ _10858_ registers\[41\]\[61\] _11585_ VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__mux2_1
XANTENNA_953 _10439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_964 _10852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_975 _11158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16432_ _14930_ _14933_ _14934_ _14935_ VGND VGND VPWR VPWR _14936_ sky130_fd_sc_hd__o211a_2
X_19220_ registers\[56\]\[24\] registers\[57\]\[24\] registers\[58\]\[24\] registers\[59\]\[24\]
+ _05958_ _05748_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__mux4_1
X_28418_ _12600_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_986 _11657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29398_ _09670_ registers\[21\]\[6\] _13140_ VGND VGND VPWR VPWR _13147_ sky130_fd_sc_hd__mux2_1
XANTENNA_997 _11818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19151_ registers\[36\]\[22\] registers\[37\]\[22\] registers\[38\]\[22\] registers\[39\]\[22\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__mux4_1
X_28349_ registers\[2\]\[52\] _10414_ _12561_ VGND VGND VPWR VPWR _12564_ sky130_fd_sc_hd__mux2_1
X_16363_ _14862_ _14868_ _14554_ _14556_ VGND VGND VPWR VPWR _14869_ sky130_fd_sc_hd__o211a_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18102_ registers\[56\]\[58\] registers\[57\]\[58\] registers\[58\]\[58\] registers\[59\]\[58\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__mux4_1
XFILLER_158_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31360_ _14134_ VGND VGND VPWR VPWR _14179_ sky130_fd_sc_hd__buf_4
X_19082_ _05755_ _05823_ _05824_ _05759_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__a22o_1
X_16294_ registers\[12\]\[6\] registers\[13\]\[6\] registers\[14\]\[6\] registers\[15\]\[6\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14802_ sky130_fd_sc_hd__mux4_1
XFILLER_201_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30311_ registers\[15\]\[55\] _13050_ _13621_ VGND VGND VPWR VPWR _13627_ sky130_fd_sc_hd__mux2_1
X_18033_ _04783_ _04790_ _04797_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__or4_4
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31291_ registers\[7\]\[7\] net62 _14135_ VGND VGND VPWR VPWR _14143_ sky130_fd_sc_hd__mux2_1
X_33030_ clknet_leaf_199_CLK _01144_ VGND VGND VPWR VPWR registers\[52\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_30242_ registers\[15\]\[22\] _12981_ _13588_ VGND VGND VPWR VPWR _13591_ sky130_fd_sc_hd__mux2_1
XFILLER_67_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30173_ _13554_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19984_ registers\[40\]\[46\] registers\[41\]\[46\] registers\[42\]\[46\] registers\[43\]\[46\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux4_1
XFILLER_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18935_ registers\[60\]\[16\] registers\[61\]\[16\] registers\[62\]\[16\] registers\[63\]\[16\]
+ _05619_ _05413_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__mux4_1
XFILLER_171_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34981_ clknet_leaf_448_CLK _03095_ VGND VGND VPWR VPWR registers\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1330 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1341 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1352 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33932_ clknet_leaf_168_CLK _02046_ VGND VGND VPWR VPWR registers\[38\]\[62\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1363 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_9_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18866_ _05078_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__buf_6
XFILLER_239_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1374 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1385 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1396 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17817_ registers\[24\]\[49\] registers\[25\]\[49\] registers\[26\]\[49\] registers\[27\]\[49\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__mux4_1
X_33863_ clknet_leaf_218_CLK _01977_ VGND VGND VPWR VPWR registers\[3\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ registers\[44\]\[12\] registers\[45\]\[12\] registers\[46\]\[12\] registers\[47\]\[12\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__mux4_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35602_ clknet_leaf_106_CLK _03716_ VGND VGND VPWR VPWR registers\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32814_ clknet_leaf_368_CLK _00928_ VGND VGND VPWR VPWR registers\[55\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_17748_ registers\[28\]\[47\] registers\[29\]\[47\] registers\[30\]\[47\] registers\[31\]\[47\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__mux4_1
X_33794_ clknet_leaf_248_CLK _01908_ VGND VGND VPWR VPWR registers\[40\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35533_ clknet_leaf_145_CLK _03647_ VGND VGND VPWR VPWR registers\[13\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_32745_ clknet_leaf_424_CLK _00859_ VGND VGND VPWR VPWR registers\[56\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_17679_ registers\[20\]\[45\] registers\[21\]\[45\] registers\[22\]\[45\] registers\[23\]\[45\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__mux4_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19418_ _06130_ _06137_ _06144_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__or4_4
X_35464_ clknet_leaf_155_CLK _03578_ VGND VGND VPWR VPWR registers\[14\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_20690_ _07388_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__buf_4
X_32676_ clknet_leaf_440_CLK _00790_ VGND VGND VPWR VPWR registers\[57\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34415_ clknet_leaf_395_CLK _02529_ VGND VGND VPWR VPWR registers\[30\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_31627_ _14319_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__clkbuf_1
X_19349_ registers\[32\]\[28\] registers\[33\]\[28\] registers\[34\]\[28\] registers\[35\]\[28\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux4_1
X_35395_ clknet_leaf_227_CLK _03509_ VGND VGND VPWR VPWR registers\[15\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22360_ _09007_ _09010_ _08740_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__o21ba_1
X_34346_ clknet_leaf_405_CLK _02460_ VGND VGND VPWR VPWR registers\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31558_ _14283_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21311_ _07328_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__clkbuf_4
X_22291_ registers\[56\]\[46\] registers\[57\]\[46\] registers\[58\]\[46\] registers\[59\]\[46\]
+ _08880_ _08670_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__mux4_1
X_30509_ _09699_ registers\[13\]\[20\] _13731_ VGND VGND VPWR VPWR _13732_ sky130_fd_sc_hd__mux2_1
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31489_ _09769_ registers\[6\]\[37\] _14239_ VGND VGND VPWR VPWR _14247_ sky130_fd_sc_hd__mux2_1
X_34277_ clknet_leaf_57_CLK _02391_ VGND VGND VPWR VPWR registers\[32\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21242_ registers\[8\]\[16\] registers\[9\]\[16\] registers\[10\]\[16\] registers\[11\]\[16\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__mux4_1
X_36016_ clknet_leaf_369_CLK _04130_ VGND VGND VPWR VPWR registers\[63\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_24030_ _10190_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__clkbuf_1
X_33228_ clknet_leaf_143_CLK _01342_ VGND VGND VPWR VPWR registers\[4\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21173_ _07648_ _07856_ _07857_ _07652_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__a22o_1
X_33159_ clknet_leaf_259_CLK _01273_ VGND VGND VPWR VPWR registers\[50\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_20124_ _06816_ _06823_ _06830_ _06837_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__or4_4
XFILLER_120_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25981_ _10835_ registers\[46\]\[50\] _11285_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__mux2_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27720_ _12221_ VGND VGND VPWR VPWR _12233_ sky130_fd_sc_hd__buf_6
X_20055_ registers\[32\]\[48\] registers\[33\]\[48\] registers\[34\]\[48\] registers\[35\]\[48\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__mux4_1
X_24932_ _10698_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27651_ registers\[34\]\[41\] _10391_ _12195_ VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__mux2_1
X_24863_ _10662_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26602_ _10781_ registers\[41\]\[24\] _11608_ VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__mux2_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23814_ _09626_ registers\[29\]\[53\] _10072_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__mux2_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ _12160_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__clkbuf_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24794_ _09588_ registers\[54\]\[35\] _10620_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__mux2_1
XANTENNA_205 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_216 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29321_ _13106_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__clkbuf_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26533_ _10848_ registers\[42\]\[56\] _11569_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__mux2_1
XFILLER_42_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23745_ _09556_ registers\[29\]\[20\] _10039_ VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__mux2_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20957_ _07324_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__clkbuf_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29252_ _13070_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__clkbuf_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26464_ _10779_ registers\[42\]\[23\] _11536_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__mux2_1
X_23676_ registers\[61\]\[53\] _09804_ _09998_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__mux2_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _07275_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__buf_4
X_28203_ _11828_ registers\[30\]\[47\] _12479_ VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__mux2_1
X_25415_ _10819_ registers\[50\]\[42\] _10981_ VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__mux2_1
X_22627_ registers\[16\]\[55\] registers\[17\]\[55\] registers\[18\]\[55\] registers\[19\]\[55\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__mux4_1
XFILLER_139_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29183_ registers\[23\]\[42\] _13023_ _13019_ VGND VGND VPWR VPWR _13024_ sky130_fd_sc_hd__mux2_1
XFILLER_41_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26395_ _11503_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28134_ _11759_ registers\[30\]\[14\] _12446_ VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__mux2_1
X_25346_ _10947_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__clkbuf_1
X_22558_ registers\[12\]\[53\] registers\[13\]\[53\] registers\[14\]\[53\] registers\[15\]\[53\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__mux4_1
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28065_ _12414_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__clkbuf_1
X_21509_ _08181_ _08184_ _08087_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__o21ba_1
XFILLER_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25277_ _10817_ registers\[51\]\[41\] _10909_ VGND VGND VPWR VPWR _10911_ sky130_fd_sc_hd__mux2_1
X_22489_ registers\[4\]\[51\] registers\[5\]\[51\] registers\[6\]\[51\] registers\[7\]\[51\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__mux4_1
XFILLER_182_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27016_ _11860_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24228_ _09632_ registers\[58\]\[56\] _10288_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__mux2_1
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1002 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24159_ _09563_ registers\[58\]\[23\] _10255_ VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16981_ registers\[44\]\[26\] registers\[45\]\[26\] registers\[46\]\[26\] registers\[47\]\[26\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15469_ sky130_fd_sc_hd__mux4_1
XFILLER_27_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28967_ registers\[24\]\[25\] _10357_ _12883_ VGND VGND VPWR VPWR _12889_ sky130_fd_sc_hd__mux2_1
XFILLER_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18720_ registers\[36\]\[10\] registers\[37\]\[10\] registers\[38\]\[10\] registers\[39\]\[10\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__mux4_1
XFILLER_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27918_ _12292_ VGND VGND VPWR VPWR _12337_ sky130_fd_sc_hd__buf_4
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28898_ _12852_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__clkbuf_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18651_ registers\[56\]\[8\] registers\[57\]\[8\] registers\[58\]\[8\] registers\[59\]\[8\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__mux4_1
X_27849_ registers\[32\]\[7\] _10319_ _12293_ VGND VGND VPWR VPWR _12301_ sky130_fd_sc_hd__mux2_1
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _15825_ _04384_ _04385_ _15828_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a22o_1
XFILLER_114_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30860_ _09817_ registers\[11\]\[59\] _13906_ VGND VGND VPWR VPWR _13916_ sky130_fd_sc_hd__mux2_1
XFILLER_91_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ registers\[60\]\[6\] registers\[61\]\[6\] registers\[62\]\[6\] registers\[63\]\[6\]
+ _05276_ _05093_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__mux4_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29519_ _12933_ _11010_ VGND VGND VPWR VPWR _13210_ sky130_fd_sc_hd__nor2_8
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ registers\[0\]\[41\] registers\[1\]\[41\] registers\[2\]\[41\] registers\[3\]\[41\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__mux4_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30791_ _09744_ registers\[11\]\[26\] _13873_ VGND VGND VPWR VPWR _13880_ sky130_fd_sc_hd__mux2_1
XFILLER_33_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_750 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_260_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_260_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_761 _07398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32530_ clknet_leaf_76_CLK _00644_ VGND VGND VPWR VPWR registers\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17464_ registers\[24\]\[39\] registers\[25\]\[39\] registers\[26\]\[39\] registers\[27\]\[39\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15939_ sky130_fd_sc_hd__mux4_1
XANTENNA_772 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_783 _08639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_794 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16415_ registers\[32\]\[10\] registers\[33\]\[10\] registers\[34\]\[10\] registers\[35\]\[10\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _14919_ sky130_fd_sc_hd__mux4_1
X_19203_ registers\[24\]\[23\] registers\[25\]\[23\] registers\[26\]\[23\] registers\[27\]\[23\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__mux4_1
XFILLER_207_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32461_ clknet_leaf_145_CLK _00575_ VGND VGND VPWR VPWR registers\[29\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_17395_ registers\[28\]\[37\] registers\[29\]\[37\] registers\[30\]\[37\] registers\[31\]\[37\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15872_ sky130_fd_sc_hd__mux4_1
X_34200_ clknet_leaf_85_CLK _02314_ VGND VGND VPWR VPWR registers\[33\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1083 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16346_ registers\[36\]\[8\] registers\[37\]\[8\] registers\[38\]\[8\] registers\[39\]\[8\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _14852_ sky130_fd_sc_hd__mux4_1
X_31412_ _09648_ registers\[6\]\[0\] _14206_ VGND VGND VPWR VPWR _14207_ sky130_fd_sc_hd__mux2_1
XFILLER_13_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19134_ registers\[16\]\[21\] registers\[17\]\[21\] registers\[18\]\[21\] registers\[19\]\[21\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__mux4_1
X_32392_ clknet_leaf_178_CLK _00506_ VGND VGND VPWR VPWR registers\[61\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_35180_ clknet_leaf_396_CLK _03294_ VGND VGND VPWR VPWR registers\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34131_ clknet_leaf_120_CLK _02245_ VGND VGND VPWR VPWR registers\[34\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_19065_ _05787_ _05794_ _05801_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__or4_1
X_31343_ _14170_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__clkbuf_1
X_16277_ _14655_ _14783_ _14784_ _14658_ VGND VGND VPWR VPWR _14785_ sky130_fd_sc_hd__a22o_1
XFILLER_173_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18016_ registers\[52\]\[55\] registers\[53\]\[55\] registers\[54\]\[55\] registers\[55\]\[55\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__mux4_1
XFILLER_103_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34062_ clknet_leaf_132_CLK _02176_ VGND VGND VPWR VPWR registers\[35\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_31274_ _14133_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_13_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_13_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_172_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30225_ registers\[15\]\[14\] _12964_ _13577_ VGND VGND VPWR VPWR _13582_ sky130_fd_sc_hd__mux2_1
X_33013_ clknet_leaf_352_CLK _01127_ VGND VGND VPWR VPWR registers\[52\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30156_ _13545_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19967_ _05053_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__buf_4
XFILLER_86_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18918_ _05496_ _05664_ _05665_ _05499_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__a22o_1
X_34964_ clknet_leaf_98_CLK _03078_ VGND VGND VPWR VPWR registers\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_28_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_28_0_CLK sky130_fd_sc_hd__clkbuf_8
X_30087_ _13509_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__clkbuf_1
X_19898_ _06441_ _06616_ _06617_ _06445_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__a22o_1
XANTENNA_1160 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1171 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1182 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33915_ clknet_leaf_282_CLK _02029_ VGND VGND VPWR VPWR registers\[38\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18849_ _05593_ _05598_ _05494_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1193 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34895_ clknet_leaf_114_CLK _03009_ VGND VGND VPWR VPWR registers\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33846_ clknet_leaf_317_CLK _01960_ VGND VGND VPWR VPWR registers\[3\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_21860_ registers\[20\]\[33\] registers\[21\]\[33\] registers\[22\]\[33\] registers\[23\]\[33\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__mux4_1
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20811_ _07440_ _07504_ _07505_ _07443_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__a22o_1
XFILLER_110_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21791_ _08423_ _08457_ _08458_ _08428_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__a22o_1
X_33777_ clknet_leaf_347_CLK _01891_ VGND VGND VPWR VPWR registers\[40\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_30989_ registers\[10\]\[56\] _13052_ _13977_ VGND VGND VPWR VPWR _13984_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_251_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_251_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23530_ _09617_ registers\[19\]\[49\] _09914_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__mux2_1
X_35516_ clknet_leaf_305_CLK _03630_ VGND VGND VPWR VPWR registers\[13\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_20742_ _07433_ _07436_ _07437_ _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__a22o_1
XFILLER_211_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32728_ clknet_leaf_67_CLK _00842_ VGND VGND VPWR VPWR registers\[56\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23461_ _09548_ registers\[19\]\[16\] _09881_ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__mux2_1
X_35447_ clknet_leaf_313_CLK _03561_ VGND VGND VPWR VPWR registers\[14\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_20673_ _07274_ VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__buf_12
X_32659_ clknet_leaf_70_CLK _00773_ VGND VGND VPWR VPWR registers\[57\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25200_ _10870_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_1
X_22412_ _08953_ _09060_ _09061_ _08956_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__a22o_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26180_ _11390_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
X_23392_ registers\[39\]\[49\] _09795_ _09840_ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__mux2_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35378_ clknet_leaf_382_CLK _03492_ VGND VGND VPWR VPWR registers\[15\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25131_ net40 VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__buf_2
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22343_ _08958_ _08993_ _08994_ _08961_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__a22o_1
X_34329_ clknet_leaf_21_CLK _02443_ VGND VGND VPWR VPWR registers\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25062_ _10778_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
X_22274_ _08924_ _08927_ _08759_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__o21ba_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24013_ _10181_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21225_ registers\[40\]\[16\] registers\[41\]\[16\] registers\[42\]\[16\] registers\[43\]\[16\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__mux4_1
X_29870_ registers\[18\]\[38\] _13014_ _13386_ VGND VGND VPWR VPWR _13395_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28821_ _12789_ VGND VGND VPWR VPWR _12812_ sky130_fd_sc_hd__buf_4
XFILLER_219_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21156_ _07838_ _07841_ _07744_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__o21ba_1
X_20107_ registers\[52\]\[49\] registers\[53\]\[49\] registers\[54\]\[49\] registers\[55\]\[49\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__mux4_1
X_28752_ _11837_ registers\[26\]\[51\] _12774_ VGND VGND VPWR VPWR _12776_ sky130_fd_sc_hd__mux2_1
X_21087_ _07753_ _07760_ _07767_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__or4_1
X_25964_ _10819_ registers\[46\]\[42\] _11274_ VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__mux2_1
XFILLER_246_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27703_ _12224_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__clkbuf_1
X_20038_ registers\[8\]\[47\] registers\[9\]\[47\] registers\[10\]\[47\] registers\[11\]\[47\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__mux4_1
X_24915_ _10689_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25895_ _11240_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
X_28683_ _12739_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__clkbuf_1
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_490_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_490_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24846_ _09640_ registers\[54\]\[60\] _10586_ VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__mux2_1
X_27634_ registers\[34\]\[33\] _10374_ _12184_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__mux2_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27565_ registers\[34\]\[0\] _10303_ _12151_ VGND VGND VPWR VPWR _12152_ sky130_fd_sc_hd__mux2_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24777_ _09571_ registers\[54\]\[27\] _10609_ VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__mux2_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21989_ registers\[4\]\[37\] registers\[5\]\[37\] registers\[6\]\[37\] registers\[7\]\[37\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__mux4_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_242_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_242_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26516_ _10831_ registers\[42\]\[48\] _11558_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__mux2_1
X_29304_ _13097_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__clkbuf_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _09540_ registers\[29\]\[12\] _10028_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__mux2_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27496_ _12114_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29235_ registers\[23\]\[59\] _13058_ _13040_ VGND VGND VPWR VPWR _13059_ sky130_fd_sc_hd__mux2_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26447_ _10762_ registers\[42\]\[15\] _11525_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__mux2_1
XFILLER_169_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23659_ registers\[61\]\[45\] _09786_ _09987_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__mux2_1
XFILLER_109_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ registers\[28\]\[3\] registers\[29\]\[3\] registers\[30\]\[3\] registers\[31\]\[3\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14711_ sky130_fd_sc_hd__mux4_1
X_17180_ registers\[0\]\[31\] registers\[1\]\[31\] registers\[2\]\[31\] registers\[3\]\[31\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15663_ sky130_fd_sc_hd__mux4_1
X_29166_ net31 VGND VGND VPWR VPWR _13012_ sky130_fd_sc_hd__clkbuf_4
X_26378_ _11494_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16131_ registers\[20\]\[1\] registers\[21\]\[1\] registers\[22\]\[1\] registers\[23\]\[1\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14644_ sky130_fd_sc_hd__mux4_1
X_28117_ _11742_ registers\[30\]\[6\] _12435_ VGND VGND VPWR VPWR _12442_ sky130_fd_sc_hd__mux2_1
XFILLER_35_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25329_ _10733_ registers\[50\]\[1\] _10937_ VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__mux2_1
X_29097_ _12965_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28048_ _12405_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__clkbuf_1
X_16062_ _14529_ VGND VGND VPWR VPWR _14576_ sky130_fd_sc_hd__buf_12
XFILLER_157_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30010_ registers\[17\]\[40\] _13018_ _13468_ VGND VGND VPWR VPWR _13469_ sky130_fd_sc_hd__mux2_1
X_19821_ registers\[44\]\[41\] registers\[45\]\[41\] registers\[46\]\[41\] registers\[47\]\[41\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__mux4_1
XFILLER_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29999_ registers\[17\]\[35\] _13008_ _13457_ VGND VGND VPWR VPWR _13463_ sky130_fd_sc_hd__mux2_1
XFILLER_68_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19752_ _06433_ _06474_ _06475_ _06439_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__a22o_1
X_16964_ _15139_ _15451_ _15452_ _15142_ VGND VGND VPWR VPWR _15453_ sky130_fd_sc_hd__a22o_1
XFILLER_46_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18703_ _05350_ _05455_ _05456_ _05353_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a22o_1
XFILLER_209_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31961_ clknet_leaf_4_CLK _00130_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
X_19683_ _06098_ _06407_ _06408_ _06102_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__a22o_1
X_16895_ registers\[0\]\[23\] registers\[1\]\[23\] registers\[2\]\[23\] registers\[3\]\[23\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15386_ sky130_fd_sc_hd__mux4_1
XFILLER_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33700_ clknet_leaf_57_CLK _01814_ VGND VGND VPWR VPWR registers\[41\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_481_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_481_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18634_ registers\[16\]\[7\] registers\[17\]\[7\] registers\[18\]\[7\] registers\[19\]\[7\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__mux4_1
X_30912_ _13943_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34680_ clknet_leaf_428_CLK _02794_ VGND VGND VPWR VPWR registers\[26\]\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31892_ _09766_ registers\[49\]\[36\] _14452_ VGND VGND VPWR VPWR _14459_ sky130_fd_sc_hd__mux2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33631_ clknet_leaf_33_CLK _01745_ VGND VGND VPWR VPWR registers\[42\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_30843_ _13907_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__clkbuf_1
X_18565_ _05137_ _05321_ _05322_ _05147_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__a22o_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_233_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_233_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17516_ _15956_ _15965_ _04288_ _04302_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__or4_1
XFILLER_221_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33562_ clknet_leaf_32_CLK _01676_ VGND VGND VPWR VPWR registers\[43\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_18496_ _05250_ _05255_ _05134_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__o21ba_1
X_30774_ _09695_ registers\[11\]\[18\] _13862_ VGND VGND VPWR VPWR _13871_ sky130_fd_sc_hd__mux2_1
XFILLER_233_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_580 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_591 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35301_ clknet_leaf_449_CLK _03415_ VGND VGND VPWR VPWR registers\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_32513_ clknet_leaf_233_CLK _00627_ VGND VGND VPWR VPWR registers\[60\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17447_ registers\[36\]\[39\] registers\[37\]\[39\] registers\[38\]\[39\] registers\[39\]\[39\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _15922_ sky130_fd_sc_hd__mux4_1
X_33493_ clknet_leaf_124_CLK _01607_ VGND VGND VPWR VPWR registers\[44\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35232_ clknet_leaf_2_CLK _03346_ VGND VGND VPWR VPWR registers\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_32444_ clknet_leaf_187_CLK _00558_ VGND VGND VPWR VPWR registers\[29\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17378_ registers\[56\]\[37\] registers\[57\]\[37\] registers\[58\]\[37\] registers\[59\]\[37\]
+ _15752_ _15542_ VGND VGND VPWR VPWR _15855_ sky130_fd_sc_hd__mux4_1
X_19117_ _05547_ _05857_ _05858_ _05550_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__a22o_1
X_16329_ registers\[12\]\[7\] registers\[13\]\[7\] registers\[14\]\[7\] registers\[15\]\[7\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14836_ sky130_fd_sc_hd__mux4_1
X_35163_ clknet_leaf_21_CLK _03277_ VGND VGND VPWR VPWR registers\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_32375_ clknet_leaf_331_CLK _00489_ VGND VGND VPWR VPWR registers\[61\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_34114_ clknet_leaf_247_CLK _02228_ VGND VGND VPWR VPWR registers\[35\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31326_ _14161_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__clkbuf_1
X_19048_ registers\[52\]\[19\] registers\[53\]\[19\] registers\[54\]\[19\] registers\[55\]\[19\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__mux4_1
XFILLER_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35094_ clknet_leaf_87_CLK _03208_ VGND VGND VPWR VPWR registers\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xoutput201 net201 VGND VGND VPWR VPWR D2[52] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR D2[62] sky130_fd_sc_hd__buf_2
XFILLER_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31257_ registers\[8\]\[55\] net51 _14119_ VGND VGND VPWR VPWR _14125_ sky130_fd_sc_hd__mux2_1
X_34045_ clknet_leaf_276_CLK _02159_ VGND VGND VPWR VPWR registers\[36\]\[47\] sky130_fd_sc_hd__dfxtp_1
Xoutput223 net223 VGND VGND VPWR VPWR D3[14] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR D3[24] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR D3[34] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR D3[44] sky130_fd_sc_hd__buf_2
XFILLER_88_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21010_ _07386_ _07698_ _07699_ _07396_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__a22o_1
Xoutput267 net267 VGND VGND VPWR VPWR D3[54] sky130_fd_sc_hd__buf_2
X_30208_ registers\[15\]\[6\] _12947_ _13566_ VGND VGND VPWR VPWR _13573_ sky130_fd_sc_hd__mux2_1
XFILLER_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput278 net278 VGND VGND VPWR VPWR D3[6] sky130_fd_sc_hd__buf_2
X_31188_ registers\[8\]\[22\] net15 _14086_ VGND VGND VPWR VPWR _14089_ sky130_fd_sc_hd__mux2_1
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30139_ _13536_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__clkbuf_1
X_35996_ clknet_leaf_55_CLK _04110_ VGND VGND VPWR VPWR registers\[63\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34947_ clknet_leaf_204_CLK _03061_ VGND VGND VPWR VPWR registers\[22\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22961_ _09569_ registers\[62\]\[26\] _09557_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__mux2_1
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24700_ _10575_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_472_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_472_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_210_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21912_ _08572_ _08575_ _08405_ _08406_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__o211a_1
X_25680_ _11126_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22892_ net45 VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__clkbuf_4
X_34878_ clknet_leaf_186_CLK _02992_ VGND VGND VPWR VPWR registers\[23\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24631_ _10539_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33829_ clknet_leaf_464_CLK _01943_ VGND VGND VPWR VPWR registers\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_21843_ registers\[60\]\[33\] registers\[61\]\[33\] registers\[62\]\[33\] registers\[63\]\[33\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__mux4_1
XFILLER_58_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_224_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_224_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27350_ _12037_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__clkbuf_1
X_24562_ _10501_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21774_ _08326_ _08440_ _08441_ _08332_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__a22o_1
XFILLER_70_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26301_ _11442_ VGND VGND VPWR VPWR _11454_ sky130_fd_sc_hd__buf_4
XFILLER_93_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23513_ _09915_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__clkbuf_1
X_27281_ _11853_ registers\[37\]\[59\] _11991_ VGND VGND VPWR VPWR _12001_ sky130_fd_sc_hd__mux2_1
X_20725_ _07355_ _07421_ _07422_ _07367_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__a22o_1
XFILLER_93_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24493_ _10465_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29020_ registers\[24\]\[50\] _10409_ _12916_ VGND VGND VPWR VPWR _12917_ sky130_fd_sc_hd__mux2_1
XFILLER_180_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26232_ _10817_ registers\[44\]\[41\] _11416_ VGND VGND VPWR VPWR _11418_ sky130_fd_sc_hd__mux2_1
XFILLER_211_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23444_ _09531_ registers\[19\]\[8\] _09870_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__mux2_1
X_20656_ _07295_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26163_ _11381_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23375_ _09841_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
X_20587_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25114_ _10813_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__clkbuf_1
X_22326_ _07356_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__buf_4
XFILLER_164_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26094_ _11300_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__buf_4
XFILLER_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29922_ registers\[18\]\[63\] _13066_ _13352_ VGND VGND VPWR VPWR _13422_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25045_ _10766_ registers\[52\]\[17\] _10752_ VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__mux2_1
XFILLER_156_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22257_ _08812_ _08909_ _08910_ _08815_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__a22o_1
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21208_ _07289_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29853_ _13352_ VGND VGND VPWR VPWR _13386_ sky130_fd_sc_hd__buf_4
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22188_ _08805_ _08842_ _08843_ _08810_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__a22o_1
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28804_ _12803_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21139_ _07648_ _07823_ _07824_ _07652_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__a22o_1
X_29784_ _13349_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__clkbuf_1
X_26996_ net52 VGND VGND VPWR VPWR _11847_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28735_ _11820_ registers\[26\]\[43\] _12763_ VGND VGND VPWR VPWR _12767_ sky130_fd_sc_hd__mux2_1
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25947_ _10802_ registers\[46\]\[34\] _11263_ VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__mux2_1
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_463_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_463_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16680_ registers\[0\]\[17\] registers\[1\]\[17\] registers\[2\]\[17\] registers\[3\]\[17\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15177_ sky130_fd_sc_hd__mux4_1
XFILLER_47_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25878_ _10733_ registers\[46\]\[1\] _11230_ VGND VGND VPWR VPWR _11232_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28666_ _11750_ registers\[26\]\[10\] _12730_ VGND VGND VPWR VPWR _12731_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24829_ _10644_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27617_ registers\[34\]\[25\] _10357_ _12173_ VGND VGND VPWR VPWR _12179_ sky130_fd_sc_hd__mux2_1
XFILLER_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28597_ _12694_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__clkbuf_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_215_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_215_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _05080_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__buf_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27548_ _12141_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__clkbuf_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _15677_ _15778_ _15779_ _15682_ VGND VGND VPWR VPWR _15780_ sky130_fd_sc_hd__a22o_1
XFILLER_214_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18281_ net78 VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__buf_6
XFILLER_163_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27479_ _12105_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29218_ _13047_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17232_ _15713_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30490_ _09681_ registers\[13\]\[11\] _13720_ VGND VGND VPWR VPWR _13722_ sky130_fd_sc_hd__mux2_1
XFILLER_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17163_ _15613_ _15622_ _15632_ _15646_ VGND VGND VPWR VPWR _15647_ sky130_fd_sc_hd__or4_4
X_29149_ registers\[23\]\[31\] _13000_ _12998_ VGND VGND VPWR VPWR _13001_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16114_ registers\[48\]\[1\] registers\[49\]\[1\] registers\[50\]\[1\] registers\[51\]\[1\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14627_ sky130_fd_sc_hd__mux4_1
X_32160_ clknet_leaf_16_CLK _00274_ VGND VGND VPWR VPWR registers\[39\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17094_ registers\[36\]\[29\] registers\[37\]\[29\] registers\[38\]\[29\] registers\[39\]\[29\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15579_ sky130_fd_sc_hd__mux4_1
X_31111_ _13992_ VGND VGND VPWR VPWR _14048_ sky130_fd_sc_hd__buf_4
X_16045_ _14502_ VGND VGND VPWR VPWR _14559_ sky130_fd_sc_hd__buf_8
X_32091_ clknet_leaf_489_CLK _00004_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dfxtp_1
XFILLER_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31042_ registers\[0\]\[17\] _12970_ _14004_ VGND VGND VPWR VPWR _14012_ sky130_fd_sc_hd__mux2_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19804_ registers\[16\]\[40\] registers\[17\]\[40\] registers\[18\]\[40\] registers\[19\]\[40\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__mux4_1
X_35850_ clknet_leaf_153_CLK _03964_ VGND VGND VPWR VPWR registers\[8\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17996_ registers\[24\]\[54\] registers\[25\]\[54\] registers\[26\]\[54\] registers\[27\]\[54\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux4_1
XFILLER_78_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34801_ clknet_leaf_384_CLK _02915_ VGND VGND VPWR VPWR registers\[24\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19735_ registers\[28\]\[38\] registers\[29\]\[38\] registers\[30\]\[38\] registers\[31\]\[38\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__mux4_1
X_35781_ clknet_leaf_228_CLK _03895_ VGND VGND VPWR VPWR registers\[0\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_16947_ registers\[32\]\[25\] registers\[33\]\[25\] registers\[34\]\[25\] registers\[35\]\[25\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15436_ sky130_fd_sc_hd__mux4_1
X_32993_ clknet_leaf_44_CLK _01107_ VGND VGND VPWR VPWR registers\[52\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_454_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_454_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_225_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34732_ clknet_leaf_410_CLK _02846_ VGND VGND VPWR VPWR registers\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31944_ _09821_ registers\[49\]\[61\] _14418_ VGND VGND VPWR VPWR _14486_ sky130_fd_sc_hd__mux2_1
X_19666_ _06389_ _06392_ _06194_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__o21ba_1
X_16878_ _15346_ _15353_ _15360_ _15369_ VGND VGND VPWR VPWR _15370_ sky130_fd_sc_hd__or4_4
XFILLER_237_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18617_ _05204_ _05369_ _05372_ _05207_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__a22o_1
XFILLER_168_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34663_ clknet_leaf_449_CLK _02777_ VGND VGND VPWR VPWR registers\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_19597_ _06300_ _06309_ _06316_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__or4_1
X_31875_ _09749_ registers\[49\]\[28\] _14441_ VGND VGND VPWR VPWR _14450_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_206_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_206_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33614_ clknet_leaf_131_CLK _01728_ VGND VGND VPWR VPWR registers\[42\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_18548_ registers\[48\]\[5\] registers\[49\]\[5\] registers\[50\]\[5\] registers\[51\]\[5\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux4_1
X_30826_ _13898_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__clkbuf_1
X_34594_ clknet_leaf_473_CLK _02708_ VGND VGND VPWR VPWR registers\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_33545_ clknet_leaf_255_CLK _01659_ VGND VGND VPWR VPWR registers\[44\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18479_ _05204_ _05237_ _05238_ _05207_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__a22o_1
XFILLER_209_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30757_ _13850_ VGND VGND VPWR VPWR _13862_ sky130_fd_sc_hd__buf_4
XFILLER_221_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20510_ registers\[20\]\[61\] registers\[21\]\[61\] registers\[22\]\[61\] registers\[23\]\[61\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__mux4_1
XFILLER_21_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33476_ clknet_leaf_251_CLK _01590_ VGND VGND VPWR VPWR registers\[45\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21490_ registers\[60\]\[23\] registers\[61\]\[23\] registers\[62\]\[23\] registers\[63\]\[23\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__mux4_1
XFILLER_18_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30688_ registers\[12\]\[41\] _13021_ _13824_ VGND VGND VPWR VPWR _13826_ sky130_fd_sc_hd__mux2_1
X_35215_ clknet_leaf_116_CLK _03329_ VGND VGND VPWR VPWR registers\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_20441_ _05040_ _07143_ _07144_ _05050_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__a22o_1
X_32427_ clknet_leaf_404_CLK _00541_ VGND VGND VPWR VPWR registers\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_36195_ clknet_leaf_28_CLK _00077_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dfxtp_1
X_35146_ clknet_leaf_153_CLK _03260_ VGND VGND VPWR VPWR registers\[1\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23160_ _09708_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__buf_4
XFILLER_147_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20372_ registers\[56\]\[57\] registers\[57\]\[57\] registers\[58\]\[57\] registers\[59\]\[57\]
+ _06987_ _06777_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__mux4_1
X_32358_ clknet_leaf_450_CLK _00472_ VGND VGND VPWR VPWR registers\[61\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22111_ registers\[20\]\[40\] registers\[21\]\[40\] registers\[22\]\[40\] registers\[23\]\[40\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__mux4_1
XFILLER_69_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31309_ _14152_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__clkbuf_1
X_23091_ registers\[39\]\[1\] _09660_ _09658_ VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__mux2_1
X_35077_ clknet_leaf_205_CLK _03191_ VGND VGND VPWR VPWR registers\[20\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32289_ clknet_leaf_479_CLK _00403_ VGND VGND VPWR VPWR registers\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22042_ _07303_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__buf_4
X_34028_ clknet_leaf_327_CLK _02142_ VGND VGND VPWR VPWR registers\[36\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26850_ net64 VGND VGND VPWR VPWR _11748_ sky130_fd_sc_hd__buf_4
XTAP_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25801_ _10791_ registers\[47\]\[29\] _11181_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26781_ _11707_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__clkbuf_1
X_35979_ clknet_leaf_150_CLK _04093_ VGND VGND VPWR VPWR registers\[6\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_23993_ _09533_ registers\[5\]\[9\] _10161_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_445_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_445_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_229_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25732_ _11153_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
X_28520_ _11740_ registers\[27\]\[5\] _12648_ VGND VGND VPWR VPWR _12654_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22944_ _09558_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28451_ _12617_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25663_ _11117_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
X_22875_ net1 VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__buf_4
XFILLER_16_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27402_ registers\[36\]\[52\] _10414_ _12062_ VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__mux2_1
X_24614_ _10530_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28382_ _12581_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__clkbuf_1
X_21826_ _07363_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__buf_4
X_25594_ _11079_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27333_ _12028_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__clkbuf_1
X_24545_ _10492_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21757_ _07392_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__buf_4
XFILLER_180_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20708_ _07356_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__clkbuf_8
X_27264_ _11992_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24476_ _10456_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
X_21688_ registers\[40\]\[29\] registers\[41\]\[29\] registers\[42\]\[29\] registers\[43\]\[29\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__mux4_1
XFILLER_106_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29003_ registers\[24\]\[42\] _10393_ _12905_ VGND VGND VPWR VPWR _12908_ sky130_fd_sc_hd__mux2_1
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26215_ _10800_ registers\[44\]\[33\] _11405_ VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__mux2_1
X_23427_ _09869_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__buf_4
XFILLER_123_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20639_ net75 VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__buf_12
X_27195_ _11767_ registers\[37\]\[18\] _11947_ VGND VGND VPWR VPWR _11956_ sky130_fd_sc_hd__mux2_1
X_26146_ _10728_ registers\[44\]\[0\] _11372_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__mux2_1
XFILLER_137_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23358_ _09832_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22309_ _08958_ _08959_ _08960_ _08961_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__a22o_1
XFILLER_124_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26077_ _11336_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23289_ net41 VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29905_ _13413_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__clkbuf_1
X_25028_ _10755_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1704 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1715 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1726 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17850_ registers\[12\]\[50\] registers\[13\]\[50\] registers\[14\]\[50\] registers\[15\]\[50\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux4_1
XANTENNA_1737 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29836_ _13377_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1748 _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1759 _07358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16801_ _14600_ VGND VGND VPWR VPWR _15295_ sky130_fd_sc_hd__clkbuf_4
XTAP_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29767_ registers\[1\]\[53\] _13046_ _13337_ VGND VGND VPWR VPWR _13341_ sky130_fd_sc_hd__mux2_1
X_17781_ _14578_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__buf_4
X_26979_ _11834_ registers\[3\]\[50\] _11835_ VGND VGND VPWR VPWR _11836_ sky130_fd_sc_hd__mux2_1
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_436_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_436_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_208_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19520_ _06036_ _06249_ _06250_ _06039_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__a22o_1
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16732_ _15224_ _15227_ _14959_ VGND VGND VPWR VPWR _15228_ sky130_fd_sc_hd__o21ba_1
X_28718_ _11803_ registers\[26\]\[35\] _12752_ VGND VGND VPWR VPWR _12758_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29698_ registers\[1\]\[20\] _12976_ _13304_ VGND VGND VPWR VPWR _13305_ sky130_fd_sc_hd__mux2_1
XFILLER_208_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19451_ registers\[16\]\[30\] registers\[17\]\[30\] registers\[18\]\[30\] registers\[19\]\[30\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__mux4_1
XFILLER_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28649_ _11734_ registers\[26\]\[2\] _12719_ VGND VGND VPWR VPWR _12722_ sky130_fd_sc_hd__mux2_1
X_16663_ registers\[40\]\[17\] registers\[41\]\[17\] registers\[42\]\[17\] registers\[43\]\[17\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15160_ sky130_fd_sc_hd__mux4_1
X_18402_ _05075_ _05106_ _05135_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__or4_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31660_ registers\[63\]\[54\] net50 _14332_ VGND VGND VPWR VPWR _14337_ sky130_fd_sc_hd__mux2_1
X_19382_ registers\[28\]\[28\] registers\[29\]\[28\] registers\[30\]\[28\] registers\[31\]\[28\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__mux4_1
XFILLER_61_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16594_ registers\[32\]\[15\] registers\[33\]\[15\] registers\[34\]\[15\] registers\[35\]\[15\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15093_ sky130_fd_sc_hd__mux4_1
XFILLER_222_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18333_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__buf_4
X_30611_ _13785_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__clkbuf_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31591_ registers\[63\]\[21\] net14 _14299_ VGND VGND VPWR VPWR _14301_ sky130_fd_sc_hd__mux2_1
XFILLER_231_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33330_ clknet_leaf_364_CLK _01444_ VGND VGND VPWR VPWR registers\[47\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_18264_ _14511_ _05026_ _05027_ _14517_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a22o_1
X_30542_ _09766_ registers\[13\]\[36\] _13742_ VGND VGND VPWR VPWR _13749_ sky130_fd_sc_hd__mux2_1
XFILLER_30_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17215_ registers\[8\]\[32\] registers\[9\]\[32\] registers\[10\]\[32\] registers\[11\]\[32\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15697_ sky130_fd_sc_hd__mux4_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33261_ clknet_leaf_379_CLK _01375_ VGND VGND VPWR VPWR registers\[48\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_18195_ registers\[60\]\[61\] registers\[61\]\[61\] registers\[62\]\[61\] registers\[63\]\[61\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux4_1
X_30473_ _09664_ registers\[13\]\[3\] _13709_ VGND VGND VPWR VPWR _13713_ sky130_fd_sc_hd__mux2_1
XFILLER_129_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35000_ clknet_leaf_309_CLK _03114_ VGND VGND VPWR VPWR registers\[21\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_32212_ clknet_leaf_287_CLK _00326_ VGND VGND VPWR VPWR registers\[9\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_17146_ _15487_ _15628_ _15629_ _15490_ VGND VGND VPWR VPWR _15630_ sky130_fd_sc_hd__a22o_1
X_33192_ clknet_leaf_401_CLK _01306_ VGND VGND VPWR VPWR registers\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32143_ clknet_leaf_133_CLK _00257_ VGND VGND VPWR VPWR registers\[39\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_17077_ _15487_ _15559_ _15562_ _15490_ VGND VGND VPWR VPWR _15563_ sky130_fd_sc_hd__a22o_1
XFILLER_143_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16028_ _14541_ VGND VGND VPWR VPWR _14542_ sky130_fd_sc_hd__buf_6
X_32074_ clknet_leaf_177_CLK _00252_ VGND VGND VPWR VPWR registers\[62\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35902_ clknet_leaf_198_CLK _04016_ VGND VGND VPWR VPWR registers\[7\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31025_ registers\[0\]\[9\] _12953_ _13993_ VGND VGND VPWR VPWR _14003_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35833_ clknet_leaf_317_CLK _03947_ VGND VGND VPWR VPWR registers\[8\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17979_ registers\[56\]\[54\] registers\[57\]\[54\] registers\[58\]\[54\] registers\[59\]\[54\]
+ _04751_ _04541_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__mux4_1
XFILLER_97_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_427_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_427_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19718_ registers\[60\]\[38\] registers\[61\]\[38\] registers\[62\]\[38\] registers\[63\]\[38\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux4_1
X_35764_ clknet_leaf_414_CLK _03878_ VGND VGND VPWR VPWR registers\[0\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_20990_ _07676_ _07679_ _07310_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__o21ba_1
X_32976_ clknet_leaf_175_CLK _01090_ VGND VGND VPWR VPWR registers\[52\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34715_ clknet_leaf_22_CLK _02829_ VGND VGND VPWR VPWR registers\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31927_ _14477_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__clkbuf_1
X_19649_ registers\[0\]\[36\] registers\[1\]\[36\] registers\[2\]\[36\] registers\[3\]\[36\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__mux4_1
X_35695_ clknet_leaf_376_CLK _03809_ VGND VGND VPWR VPWR registers\[10\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22660_ registers\[20\]\[56\] registers\[21\]\[56\] registers\[22\]\[56\] registers\[23\]\[56\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__mux4_1
X_34646_ clknet_leaf_89_CLK _02760_ VGND VGND VPWR VPWR registers\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31858_ _14418_ VGND VGND VPWR VPWR _14441_ sky130_fd_sc_hd__buf_4
XFILLER_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21611_ registers\[20\]\[26\] registers\[21\]\[26\] registers\[22\]\[26\] registers\[23\]\[26\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__mux4_1
XFILLER_55_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30809_ _13889_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__clkbuf_1
X_34577_ clknet_leaf_111_CLK _02691_ VGND VGND VPWR VPWR registers\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_22591_ registers\[4\]\[54\] registers\[5\]\[54\] registers\[6\]\[54\] registers\[7\]\[54\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31789_ registers\[59\]\[51\] net47 _14403_ VGND VGND VPWR VPWR _14405_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24330_ registers\[57\]\[27\] _10361_ _10347_ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__mux2_1
XFILLER_205_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33528_ clknet_leaf_339_CLK _01642_ VGND VGND VPWR VPWR registers\[44\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_21542_ _08080_ _08215_ _08216_ _08085_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__a22o_1
XFILLER_221_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24261_ net56 VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__buf_4
XFILLER_18_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21473_ _07388_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__clkbuf_4
X_33459_ clknet_leaf_347_CLK _01573_ VGND VGND VPWR VPWR registers\[45\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_26000_ _11295_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_51__f_CLK clknet_5_25_0_CLK VGND VGND VPWR VPWR clknet_6_51__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23212_ _09737_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__clkbuf_1
X_20424_ _07128_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__buf_4
X_36178_ clknet_leaf_92_CLK _00108_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dfxtp_1
X_24192_ _09596_ registers\[58\]\[39\] _10266_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__mux2_1
XFILLER_105_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35129_ clknet_leaf_302_CLK _03243_ VGND VGND VPWR VPWR registers\[1\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_23143_ registers\[39\]\[18\] _09695_ _09679_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__mux2_1
XFILLER_107_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20355_ _07058_ _07061_ _06866_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__o21ba_1
XFILLER_105_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27951_ _12354_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__clkbuf_1
X_23074_ net60 VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__buf_2
XTAP_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20286_ _06990_ _06994_ _06855_ _06856_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__o211a_1
XTAP_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26902_ _11783_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22025_ _08610_ _08684_ _08685_ _08613_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__a22o_1
XTAP_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27882_ _12318_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29621_ registers\[20\]\[48\] _13035_ _13255_ VGND VGND VPWR VPWR _13264_ sky130_fd_sc_hd__mux2_1
XFILLER_248_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26833_ _11736_ registers\[3\]\[3\] _11730_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__mux2_1
XFILLER_248_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_418_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_418_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29552_ registers\[20\]\[15\] _12966_ _13222_ VGND VGND VPWR VPWR _13228_ sky130_fd_sc_hd__mux2_1
X_23976_ _10162_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26764_ _11698_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__clkbuf_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28503_ _12644_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__clkbuf_1
X_25715_ registers\[48\]\[53\] _10416_ _11141_ VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__mux2_1
X_22927_ _09546_ registers\[62\]\[15\] _09536_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__mux2_1
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26695_ _11662_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__clkbuf_1
X_29483_ _13191_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28434_ _12608_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22858_ _09490_ _09493_ _07338_ _07340_ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__o211a_1
XFILLER_186_1287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25646_ registers\[48\]\[20\] _10346_ _11108_ VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__mux2_1
XFILLER_231_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21809_ registers\[48\]\[32\] registers\[49\]\[32\] registers\[50\]\[32\] registers\[51\]\[32\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__mux4_1
X_28365_ registers\[2\]\[60\] _10430_ _12505_ VGND VGND VPWR VPWR _12572_ sky130_fd_sc_hd__mux2_1
X_25577_ registers\[4\]\[53\] _10416_ _11067_ VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__mux2_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22789_ registers\[36\]\[61\] registers\[37\]\[61\] registers\[38\]\[61\] registers\[39\]\[61\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__mux4_1
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27316_ registers\[36\]\[11\] _10328_ _12018_ VGND VGND VPWR VPWR _12020_ sky130_fd_sc_hd__mux2_1
X_24528_ _10483_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28296_ registers\[2\]\[27\] _10361_ _12528_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__mux2_1
XFILLER_196_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24459_ _10447_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
X_27247_ _11983_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17000_ registers\[12\]\[26\] registers\[13\]\[26\] registers\[14\]\[26\] registers\[15\]\[26\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15488_ sky130_fd_sc_hd__mux4_1
XFILLER_184_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27178_ _11935_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_8 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26129_ _11363_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18951_ _05692_ _05697_ _05494_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1501 _07338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17902_ _14493_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__buf_8
XANTENNA_1512 _07547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1523 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18882_ _05111_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__buf_6
XTAP_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1534 _09535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1545 _10332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1556 _11513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17833_ _04340_ _04608_ _04609_ _04343_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__a22o_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29819_ _13368_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1567 _12363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1578 _13708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1589 _14510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_409_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_409_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32830_ clknet_leaf_292_CLK _00944_ VGND VGND VPWR VPWR registers\[55\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17764_ _14541_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__buf_4
XFILLER_130_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19503_ registers\[44\]\[32\] registers\[45\]\[32\] registers\[46\]\[32\] registers\[47\]\[32\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16715_ _15206_ _15208_ _15209_ _15210_ VGND VGND VPWR VPWR _15211_ sky130_fd_sc_hd__a22o_1
X_32761_ clknet_leaf_333_CLK _00875_ VGND VGND VPWR VPWR registers\[56\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17695_ _14546_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__buf_4
XFILLER_63_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34500_ clknet_leaf_224_CLK _02614_ VGND VGND VPWR VPWR registers\[2\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_19434_ registers\[52\]\[30\] registers\[53\]\[30\] registers\[54\]\[30\] registers\[55\]\[30\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__mux4_1
XFILLER_63_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31712_ _14364_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16646_ _14510_ VGND VGND VPWR VPWR _15144_ sky130_fd_sc_hd__clkbuf_4
X_35480_ clknet_leaf_444_CLK _03594_ VGND VGND VPWR VPWR registers\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_32692_ clknet_leaf_351_CLK _00806_ VGND VGND VPWR VPWR registers\[57\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34431_ clknet_leaf_306_CLK _02545_ VGND VGND VPWR VPWR registers\[30\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31643_ registers\[63\]\[46\] net41 _14321_ VGND VGND VPWR VPWR _14328_ sky130_fd_sc_hd__mux2_1
X_19365_ registers\[60\]\[28\] registers\[61\]\[28\] registers\[62\]\[28\] registers\[63\]\[28\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__mux4_1
X_16577_ _14796_ _15075_ _15076_ _14799_ VGND VGND VPWR VPWR _15077_ sky130_fd_sc_hd__a22o_1
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18316_ _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__buf_12
XFILLER_163_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34362_ clknet_leaf_60_CLK _02476_ VGND VGND VPWR VPWR registers\[31\]\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31574_ registers\[63\]\[13\] net5 _14288_ VGND VGND VPWR VPWR _14292_ sky130_fd_sc_hd__mux2_1
X_19296_ registers\[0\]\[26\] registers\[1\]\[26\] registers\[2\]\[26\] registers\[3\]\[26\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__mux4_1
XFILLER_206_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36101_ clknet_leaf_264_CLK _04215_ VGND VGND VPWR VPWR registers\[59\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33313_ clknet_leaf_34_CLK _01427_ VGND VGND VPWR VPWR registers\[47\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18247_ _14528_ _05009_ _05010_ _14537_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a22o_1
X_30525_ _09749_ registers\[13\]\[28\] _13731_ VGND VGND VPWR VPWR _13740_ sky130_fd_sc_hd__mux2_1
X_34293_ clknet_leaf_343_CLK _02407_ VGND VGND VPWR VPWR registers\[32\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_36032_ clknet_leaf_266_CLK _04146_ VGND VGND VPWR VPWR registers\[63\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_33244_ clknet_leaf_39_CLK _01358_ VGND VGND VPWR VPWR registers\[48\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_18178_ _14558_ _04943_ _04944_ _14568_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__a22o_1
X_30456_ _13703_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17129_ _15606_ _15611_ _15612_ VGND VGND VPWR VPWR _15613_ sky130_fd_sc_hd__o21ba_1
X_33175_ clknet_leaf_82_CLK _01289_ VGND VGND VPWR VPWR registers\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30387_ _13667_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__clkbuf_1
X_20140_ registers\[52\]\[50\] registers\[53\]\[50\] registers\[54\]\[50\] registers\[55\]\[50\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32126_ clknet_leaf_397_CLK _00042_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20071_ registers\[60\]\[48\] registers\[61\]\[48\] registers\[62\]\[48\] registers\[63\]\[48\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux4_1
X_32057_ clknet_leaf_332_CLK _00235_ VGND VGND VPWR VPWR registers\[62\]\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31008_ _13994_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__clkbuf_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23830_ _09642_ registers\[29\]\[61\] _10016_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__mux2_1
XFILLER_57_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35816_ clknet_leaf_460_CLK _03930_ VGND VGND VPWR VPWR registers\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35747_ clknet_leaf_464_CLK _03861_ VGND VGND VPWR VPWR registers\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_23761_ _09573_ registers\[29\]\[28\] _10039_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__mux2_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_409 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32959_ clknet_leaf_290_CLK _01073_ VGND VGND VPWR VPWR registers\[53\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_20973_ registers\[24\]\[8\] registers\[25\]\[8\] registers\[26\]\[8\] registers\[27\]\[8\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__mux4_1
X_22712_ registers\[12\]\[58\] registers\[13\]\[58\] registers\[14\]\[58\] registers\[15\]\[58\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__mux4_1
X_25500_ _11030_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26480_ _11548_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__clkbuf_1
X_23692_ registers\[61\]\[61\] _09821_ _09942_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__mux2_1
X_35678_ clknet_leaf_489_CLK _03792_ VGND VGND VPWR VPWR registers\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25431_ _10936_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__buf_6
X_34629_ clknet_leaf_219_CLK _02743_ VGND VGND VPWR VPWR registers\[27\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_22643_ registers\[48\]\[56\] registers\[49\]\[56\] registers\[50\]\[56\] registers\[51\]\[56\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__mux4_1
XFILLER_81_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25362_ _10766_ registers\[50\]\[17\] _10948_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__mux2_1
X_28150_ _12459_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__clkbuf_1
X_22574_ registers\[44\]\[54\] registers\[45\]\[54\] registers\[46\]\[54\] registers\[47\]\[54\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27101_ _11906_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_1
X_24313_ _10350_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
X_28081_ _11841_ registers\[31\]\[53\] _12419_ VGND VGND VPWR VPWR _12423_ sky130_fd_sc_hd__mux2_1
XFILLER_142_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21525_ registers\[52\]\[24\] registers\[53\]\[24\] registers\[54\]\[24\] registers\[55\]\[24\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__mux4_1
X_25293_ _10833_ registers\[51\]\[49\] _10909_ VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27032_ _11870_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__clkbuf_1
X_24244_ net1 VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__buf_4
XFILLER_120_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21456_ registers\[48\]\[22\] registers\[49\]\[22\] registers\[50\]\[22\] registers\[51\]\[22\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__mux4_1
XFILLER_108_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20407_ _05149_ _07110_ _07111_ _05159_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__a22o_1
X_24175_ _10267_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21387_ _07347_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__buf_6
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23126_ _09684_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
X_20338_ registers\[44\]\[56\] registers\[45\]\[56\] registers\[46\]\[56\] registers\[47\]\[56\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__mux4_1
XFILLER_123_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28983_ _12897_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__clkbuf_1
XTAP_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23057_ _09634_ registers\[62\]\[57\] _09620_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__mux2_1
X_27934_ _12345_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20269_ _06955_ _06962_ _06971_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__or4_4
XTAP_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22008_ _07312_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__clkbuf_4
XTAP_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27865_ _12309_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__clkbuf_1
XTAP_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29604_ _13210_ VGND VGND VPWR VPWR _13255_ sky130_fd_sc_hd__buf_4
X_26816_ _11725_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__clkbuf_1
XTAP_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27796_ registers\[33\]\[46\] _10401_ _12266_ VGND VGND VPWR VPWR _12273_ sky130_fd_sc_hd__mux2_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29535_ registers\[20\]\[7\] _12949_ _13211_ VGND VGND VPWR VPWR _13219_ sky130_fd_sc_hd__mux2_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26747_ _11689_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_1
X_23959_ _10152_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_910 _09691_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_921 _09780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16500_ _14998_ _14999_ _15000_ _15001_ VGND VGND VPWR VPWR _15002_ sky130_fd_sc_hd__a22o_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29466_ _13182_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_932 _10016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17480_ _15684_ _15952_ _15953_ _15687_ VGND VGND VPWR VPWR _15954_ sky130_fd_sc_hd__a22o_1
X_26678_ _11652_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_943 _10336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_954 _10495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_965 _10864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28417_ _11771_ registers\[28\]\[20\] _12599_ VGND VGND VPWR VPWR _12600_ sky130_fd_sc_hd__mux2_1
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16431_ _14555_ VGND VGND VPWR VPWR _14935_ sky130_fd_sc_hd__clkbuf_4
X_25629_ registers\[48\]\[12\] _10330_ _11097_ VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__mux2_1
XANTENNA_976 _11229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29397_ _13146_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_987 _11729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_998 _11818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19150_ registers\[44\]\[22\] registers\[45\]\[22\] registers\[46\]\[22\] registers\[47\]\[22\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__mux4_1
X_28348_ _12563_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16362_ _14863_ _14865_ _14866_ _14867_ VGND VGND VPWR VPWR _14868_ sky130_fd_sc_hd__a22o_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18101_ _04866_ _04869_ _04611_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__o21ba_2
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16293_ _14510_ VGND VGND VPWR VPWR _14801_ sky130_fd_sc_hd__buf_4
XFILLER_40_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19081_ registers\[52\]\[20\] registers\[53\]\[20\] registers\[54\]\[20\] registers\[55\]\[20\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__mux4_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28279_ registers\[2\]\[19\] _10344_ _12517_ VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__mux2_1
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30310_ _13626_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__clkbuf_1
X_18032_ _04800_ _04803_ _04644_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__o21ba_1
X_31290_ _14142_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30241_ _13590_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30172_ registers\[16\]\[53\] _13046_ _13550_ VGND VGND VPWR VPWR _13554_ sky130_fd_sc_hd__mux2_1
XFILLER_207_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19983_ _06700_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18934_ _05404_ _05679_ _05680_ _05410_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a22o_1
X_34980_ clknet_leaf_471_CLK _03094_ VGND VGND VPWR VPWR registers\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1320 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1331 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33931_ clknet_leaf_165_CLK _02045_ VGND VGND VPWR VPWR registers\[38\]\[61\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1342 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18865_ _05610_ _05613_ _05475_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1353 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1364 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1375 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1386 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17816_ _04590_ _04593_ _15974_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__o21ba_1
X_33862_ clknet_leaf_218_CLK _01976_ VGND VGND VPWR VPWR registers\[3\]\[56\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1397 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18796_ _05088_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__clkbuf_4
XTAP_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35601_ clknet_leaf_109_CLK _03715_ VGND VGND VPWR VPWR registers\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_32813_ clknet_leaf_374_CLK _00927_ VGND VGND VPWR VPWR registers\[55\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_17747_ _04289_ _04525_ _04526_ _04292_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__a22o_1
X_33793_ clknet_leaf_272_CLK _01907_ VGND VGND VPWR VPWR registers\[40\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35532_ clknet_leaf_150_CLK _03646_ VGND VGND VPWR VPWR registers\[13\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32744_ clknet_leaf_436_CLK _00858_ VGND VGND VPWR VPWR registers\[56\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17678_ registers\[28\]\[45\] registers\[29\]\[45\] registers\[30\]\[45\] registers\[31\]\[45\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__mux4_1
XFILLER_74_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19417_ _06147_ _06150_ _05851_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__o21ba_1
X_35463_ clknet_leaf_215_CLK _03577_ VGND VGND VPWR VPWR registers\[14\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16629_ registers\[36\]\[16\] registers\[37\]\[16\] registers\[38\]\[16\] registers\[39\]\[16\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _15127_ sky130_fd_sc_hd__mux4_1
X_32675_ clknet_leaf_441_CLK _00789_ VGND VGND VPWR VPWR registers\[57\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_34414_ clknet_leaf_387_CLK _02528_ VGND VGND VPWR VPWR registers\[30\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31626_ registers\[63\]\[38\] net32 _14310_ VGND VGND VPWR VPWR _14319_ sky130_fd_sc_hd__mux2_1
X_19348_ registers\[40\]\[28\] registers\[41\]\[28\] registers\[42\]\[28\] registers\[43\]\[28\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__mux4_1
X_35394_ clknet_leaf_239_CLK _03508_ VGND VGND VPWR VPWR registers\[15\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34345_ clknet_leaf_401_CLK _02459_ VGND VGND VPWR VPWR registers\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31557_ registers\[63\]\[5\] net56 _14277_ VGND VGND VPWR VPWR _14283_ sky130_fd_sc_hd__mux2_1
X_19279_ registers\[32\]\[26\] registers\[33\]\[26\] registers\[34\]\[26\] registers\[35\]\[26\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__mux4_1
XFILLER_206_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21310_ _07324_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__clkbuf_4
X_30508_ _13708_ VGND VGND VPWR VPWR _13731_ sky130_fd_sc_hd__buf_4
XFILLER_248_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22290_ _08939_ _08942_ _08740_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__o21ba_1
X_34276_ clknet_leaf_433_CLK _02390_ VGND VGND VPWR VPWR registers\[32\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31488_ _14246_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36015_ clknet_leaf_369_CLK _04129_ VGND VGND VPWR VPWR registers\[63\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33227_ clknet_leaf_158_CLK _01341_ VGND VGND VPWR VPWR registers\[4\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_21241_ _07275_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__buf_4
X_30439_ _09800_ registers\[14\]\[51\] _13693_ VGND VGND VPWR VPWR _13695_ sky130_fd_sc_hd__mux2_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33158_ clknet_leaf_262_CLK _01272_ VGND VGND VPWR VPWR registers\[50\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21172_ registers\[52\]\[14\] registers\[53\]\[14\] registers\[54\]\[14\] registers\[55\]\[14\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20123_ _06833_ _06836_ _06537_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32109_ clknet_leaf_468_CLK _00024_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dfxtp_1
X_25980_ _11229_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__buf_4
X_33089_ clknet_leaf_270_CLK _01203_ VGND VGND VPWR VPWR registers\[51\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20054_ registers\[40\]\[48\] registers\[41\]\[48\] registers\[42\]\[48\] registers\[43\]\[48\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__mux4_1
X_24931_ _09590_ registers\[53\]\[36\] _10691_ VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__mux2_1
XFILLER_219_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27650_ _12196_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__clkbuf_1
X_24862_ _09521_ registers\[53\]\[3\] _10658_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__mux2_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26601_ _11612_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23813_ _10075_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__clkbuf_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27581_ registers\[34\]\[8\] _10321_ _12151_ VGND VGND VPWR VPWR _12160_ sky130_fd_sc_hd__mux2_1
XFILLER_172_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24793_ _10625_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__clkbuf_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29320_ _09760_ registers\[22\]\[33\] _13102_ VGND VGND VPWR VPWR _13106_ sky130_fd_sc_hd__mux2_1
XANTENNA_217 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26532_ _11575_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_228 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23744_ _10016_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__buf_4
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _07640_ _07642_ _07645_ _07646_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__a22o_1
XANTENNA_239 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29251_ _09648_ registers\[22\]\[0\] _13069_ VGND VGND VPWR VPWR _13070_ sky130_fd_sc_hd__mux2_1
XFILLER_41_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _10001_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26463_ _11539_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20887_ _07574_ _07579_ _07339_ _07341_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__o211a_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28202_ _12486_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22626_ registers\[24\]\[55\] registers\[25\]\[55\] registers\[26\]\[55\] registers\[27\]\[55\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__mux4_1
X_25414_ _10983_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__clkbuf_1
X_26394_ _10844_ registers\[43\]\[54\] _11498_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__mux2_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29182_ net37 VGND VGND VPWR VPWR _13023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_70_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25345_ _10749_ registers\[50\]\[9\] _10937_ VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__mux2_1
X_28133_ _12450_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__clkbuf_1
X_22557_ _07305_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__buf_4
XFILLER_210_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21508_ _08080_ _08182_ _08183_ _08085_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__a22o_1
XFILLER_154_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28064_ _11824_ registers\[31\]\[45\] _12408_ VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__mux2_1
X_25276_ _10910_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22488_ registers\[12\]\[51\] registers\[13\]\[51\] registers\[14\]\[51\] registers\[15\]\[51\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__mux4_1
XFILLER_33_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27015_ _11859_ registers\[3\]\[62\] _11729_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__mux2_1
X_24227_ _10294_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21439_ _08113_ _08116_ _08087_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__o21ba_1
XFILLER_182_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24158_ _10258_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23109_ registers\[39\]\[7\] _09672_ _09658_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__mux2_1
X_24089_ _10221_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
X_28966_ _12888_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__clkbuf_1
X_16980_ _15334_ _15466_ _15467_ _15339_ VGND VGND VPWR VPWR _15468_ sky130_fd_sc_hd__a22o_1
XFILLER_122_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27917_ _12336_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__clkbuf_1
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28897_ _11847_ registers\[25\]\[56\] _12845_ VGND VGND VPWR VPWR _12852_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _05080_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__buf_4
X_27848_ _12300_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__clkbuf_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ registers\[0\]\[43\] registers\[1\]\[43\] registers\[2\]\[43\] registers\[3\]\[43\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__mux4_1
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _05077_ _05336_ _05337_ _05086_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a22o_1
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27779_ registers\[33\]\[38\] _10384_ _12255_ VGND VGND VPWR VPWR _12264_ sky130_fd_sc_hd__mux2_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29518_ _13209_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17532_ registers\[8\]\[41\] registers\[9\]\[41\] registers\[10\]\[41\] registers\[11\]\[41\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__mux4_1
XFILLER_166_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30790_ _13879_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_740 _07359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_751 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_762 _07401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29449_ _09753_ registers\[21\]\[30\] _13173_ VGND VGND VPWR VPWR _13174_ sky130_fd_sc_hd__mux2_1
X_17463_ _15934_ _15937_ _15631_ VGND VGND VPWR VPWR _15938_ sky130_fd_sc_hd__o21ba_1
XANTENNA_773 _08013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_784 _08709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_795 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19202_ _05936_ _05941_ _05837_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o21ba_1
X_16414_ registers\[40\]\[10\] registers\[41\]\[10\] registers\[42\]\[10\] registers\[43\]\[10\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14918_ sky130_fd_sc_hd__mux4_1
X_32460_ clknet_leaf_141_CLK _00574_ VGND VGND VPWR VPWR registers\[29\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_17394_ _15633_ _15869_ _15870_ _15636_ VGND VGND VPWR VPWR _15871_ sky130_fd_sc_hd__a22o_1
XFILLER_220_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31411_ _14205_ VGND VGND VPWR VPWR _14206_ sky130_fd_sc_hd__buf_4
X_19133_ registers\[24\]\[21\] registers\[25\]\[21\] registers\[26\]\[21\] registers\[27\]\[21\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__mux4_1
X_16345_ registers\[44\]\[8\] registers\[45\]\[8\] registers\[46\]\[8\] registers\[47\]\[8\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14851_ sky130_fd_sc_hd__mux4_1
XFILLER_201_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32391_ clknet_leaf_207_CLK _00505_ VGND VGND VPWR VPWR registers\[61\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34130_ clknet_leaf_122_CLK _02244_ VGND VGND VPWR VPWR registers\[34\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19064_ _05804_ _05807_ _05508_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__o21ba_1
X_31342_ registers\[7\]\[31\] net25 _14168_ VGND VGND VPWR VPWR _14170_ sky130_fd_sc_hd__mux2_1
X_16276_ registers\[36\]\[6\] registers\[37\]\[6\] registers\[38\]\[6\] registers\[39\]\[6\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14784_ sky130_fd_sc_hd__mux4_1
XFILLER_51_1371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18015_ registers\[60\]\[55\] registers\[61\]\[55\] registers\[62\]\[55\] registers\[63\]\[55\]
+ _04755_ _04549_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__mux4_1
XFILLER_173_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34061_ clknet_leaf_171_CLK _02175_ VGND VGND VPWR VPWR registers\[36\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31273_ registers\[8\]\[63\] net60 _14063_ VGND VGND VPWR VPWR _14133_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33012_ clknet_leaf_351_CLK _01126_ VGND VGND VPWR VPWR registers\[52\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30224_ _13581_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19966_ _05051_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__buf_6
X_30155_ registers\[16\]\[45\] _13029_ _13539_ VGND VGND VPWR VPWR _13545_ sky130_fd_sc_hd__mux2_1
XFILLER_113_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18917_ registers\[16\]\[15\] registers\[17\]\[15\] registers\[18\]\[15\] registers\[19\]\[15\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__mux4_1
X_34963_ clknet_leaf_97_CLK _03077_ VGND VGND VPWR VPWR registers\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19897_ registers\[52\]\[43\] registers\[53\]\[43\] registers\[54\]\[43\] registers\[55\]\[43\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__mux4_1
XANTENNA_1150 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30086_ registers\[16\]\[12\] _12960_ _13506_ VGND VGND VPWR VPWR _13509_ sky130_fd_sc_hd__mux2_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1161 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1172 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33914_ clknet_leaf_281_CLK _02028_ VGND VGND VPWR VPWR registers\[38\]\[44\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1183 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18848_ _05350_ _05596_ _05597_ _05353_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__a22o_1
X_34894_ clknet_leaf_115_CLK _03008_ VGND VGND VPWR VPWR registers\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1194 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33845_ clknet_leaf_415_CLK _01959_ VGND VGND VPWR VPWR registers\[3\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18779_ _05527_ _05530_ _05494_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__o21ba_1
X_20810_ registers\[36\]\[4\] registers\[37\]\[4\] registers\[38\]\[4\] registers\[39\]\[4\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__mux4_1
XFILLER_209_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21790_ registers\[20\]\[31\] registers\[21\]\[31\] registers\[22\]\[31\] registers\[23\]\[31\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__mux4_1
X_33776_ clknet_leaf_347_CLK _01890_ VGND VGND VPWR VPWR registers\[40\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30988_ _13983_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35515_ clknet_leaf_305_CLK _03629_ VGND VGND VPWR VPWR registers\[13\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_32727_ clknet_leaf_65_CLK _00841_ VGND VGND VPWR VPWR registers\[56\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_20741_ _07352_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__buf_4
XFILLER_180_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23460_ _09887_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
X_35446_ clknet_leaf_320_CLK _03560_ VGND VGND VPWR VPWR registers\[14\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20672_ _07354_ _07368_ _07370_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__o21ba_1
X_32658_ clknet_leaf_74_CLK _00772_ VGND VGND VPWR VPWR registers\[57\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22411_ registers\[0\]\[49\] registers\[1\]\[49\] registers\[2\]\[49\] registers\[3\]\[49\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__mux4_1
XFILLER_149_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31609_ _14276_ VGND VGND VPWR VPWR _14310_ sky130_fd_sc_hd__buf_4
X_23391_ _09849_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
X_35377_ clknet_leaf_381_CLK _03491_ VGND VGND VPWR VPWR registers\[15\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_32589_ clknet_leaf_145_CLK _00703_ VGND VGND VPWR VPWR registers\[5\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25130_ _10824_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22342_ registers\[4\]\[47\] registers\[5\]\[47\] registers\[6\]\[47\] registers\[7\]\[47\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__mux4_1
X_34328_ clknet_leaf_19_CLK _02442_ VGND VGND VPWR VPWR registers\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25061_ _10777_ registers\[52\]\[22\] _10773_ VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__mux2_1
X_34259_ clknet_leaf_120_CLK _02373_ VGND VGND VPWR VPWR registers\[32\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22273_ _08615_ _08925_ _08926_ _08618_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__a22o_1
XFILLER_219_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24012_ _09552_ registers\[5\]\[18\] _10172_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__mux2_1
XFILLER_163_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21224_ _07907_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28820_ _12811_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21155_ _07737_ _07839_ _07840_ _07742_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__a22o_1
XFILLER_104_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20106_ registers\[60\]\[49\] registers\[61\]\[49\] registers\[62\]\[49\] registers\[63\]\[49\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__mux4_1
X_28751_ _12775_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25963_ _11276_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21086_ _07770_ _07773_ _07744_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__o21ba_1
XFILLER_219_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27702_ registers\[33\]\[1\] _10307_ _12222_ VGND VGND VPWR VPWR _12224_ sky130_fd_sc_hd__mux2_1
X_20037_ _06749_ _06752_ _06512_ _06513_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__o211a_1
X_24914_ _09573_ registers\[53\]\[28\] _10680_ VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__mux2_1
X_28682_ _11767_ registers\[26\]\[18\] _12730_ VGND VGND VPWR VPWR _12739_ sky130_fd_sc_hd__mux2_1
XFILLER_74_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25894_ _10749_ registers\[46\]\[9\] _11230_ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__mux2_1
XFILLER_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27633_ _12187_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24845_ _10652_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27564_ _12150_ VGND VGND VPWR VPWR _12151_ sky130_fd_sc_hd__buf_6
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ registers\[12\]\[37\] registers\[13\]\[37\] registers\[14\]\[37\] registers\[15\]\[37\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__mux4_1
X_24776_ _10616_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29303_ _09742_ registers\[22\]\[25\] _13091_ VGND VGND VPWR VPWR _13097_ sky130_fd_sc_hd__mux2_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26515_ _11566_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _07627_ _07630_ _07399_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o21ba_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23727_ _10030_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27495_ _11797_ registers\[35\]\[32\] _12111_ VGND VGND VPWR VPWR _12114_ sky130_fd_sc_hd__mux2_1
XFILLER_215_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29234_ net55 VGND VGND VPWR VPWR _13058_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26446_ _11530_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__clkbuf_1
X_23658_ _09992_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22609_ registers\[36\]\[55\] registers\[37\]\[55\] registers\[38\]\[55\] registers\[39\]\[55\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__mux4_1
XFILLER_168_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29165_ _13011_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__clkbuf_1
X_26377_ _10827_ registers\[43\]\[46\] _11487_ VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__mux2_1
X_23589_ _09956_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16130_ registers\[28\]\[1\] registers\[29\]\[1\] registers\[30\]\[1\] registers\[31\]\[1\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _14643_ sky130_fd_sc_hd__mux4_1
X_28116_ _12441_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__clkbuf_1
X_25328_ _10938_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29096_ registers\[23\]\[14\] _12964_ _12956_ VGND VGND VPWR VPWR _12965_ sky130_fd_sc_hd__mux2_1
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16061_ registers\[12\]\[0\] registers\[13\]\[0\] registers\[14\]\[0\] registers\[15\]\[0\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _14575_ sky130_fd_sc_hd__mux4_1
XFILLER_143_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28047_ _11807_ registers\[31\]\[37\] _12397_ VGND VGND VPWR VPWR _12405_ sky130_fd_sc_hd__mux2_1
X_25259_ _10901_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19820_ _06226_ _06540_ _06541_ _06231_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__a22o_1
XFILLER_233_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29998_ _13462_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19751_ registers\[48\]\[39\] registers\[49\]\[39\] registers\[50\]\[39\] registers\[51\]\[39\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__mux4_1
X_16963_ registers\[0\]\[25\] registers\[1\]\[25\] registers\[2\]\[25\] registers\[3\]\[25\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15452_ sky130_fd_sc_hd__mux4_1
X_28949_ _12879_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18702_ registers\[4\]\[9\] registers\[5\]\[9\] registers\[6\]\[9\] registers\[7\]\[9\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__mux4_1
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_28__f_CLK clknet_5_14_0_CLK VGND VGND VPWR VPWR clknet_6_28__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31960_ clknet_leaf_4_CLK _00129_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
X_19682_ registers\[52\]\[37\] registers\[53\]\[37\] registers\[54\]\[37\] registers\[55\]\[37\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__mux4_1
X_16894_ registers\[8\]\[23\] registers\[9\]\[23\] registers\[10\]\[23\] registers\[11\]\[23\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15385_ sky130_fd_sc_hd__mux4_1
X_18633_ registers\[24\]\[7\] registers\[25\]\[7\] registers\[26\]\[7\] registers\[27\]\[7\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__mux4_1
X_30911_ registers\[10\]\[19\] _12974_ _13933_ VGND VGND VPWR VPWR _13943_ sky130_fd_sc_hd__mux2_1
XFILLER_225_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31891_ _14458_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33630_ clknet_leaf_27_CLK _01744_ VGND VGND VPWR VPWR registers\[42\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30842_ _09797_ registers\[11\]\[50\] _13906_ VGND VGND VPWR VPWR _13907_ sky130_fd_sc_hd__mux2_1
X_18564_ registers\[16\]\[5\] registers\[17\]\[5\] registers\[18\]\[5\] registers\[19\]\[5\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__mux4_1
XFILLER_40_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _04293_ _04300_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__o21ba_1
X_33561_ clknet_leaf_90_CLK _01675_ VGND VGND VPWR VPWR registers\[43\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18495_ _05119_ _05253_ _05254_ _05131_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a22o_1
X_30773_ _13870_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_570 _04863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35300_ clknet_leaf_447_CLK _03414_ VGND VGND VPWR VPWR registers\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32512_ clknet_leaf_294_CLK _00626_ VGND VGND VPWR VPWR registers\[60\]\[50\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_581 _05051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_592 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17446_ registers\[44\]\[39\] registers\[45\]\[39\] registers\[46\]\[39\] registers\[47\]\[39\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15921_ sky130_fd_sc_hd__mux4_1
X_33492_ clknet_leaf_125_CLK _01606_ VGND VGND VPWR VPWR registers\[44\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35231_ clknet_leaf_2_CLK _03345_ VGND VGND VPWR VPWR registers\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_32443_ clknet_leaf_183_CLK _00557_ VGND VGND VPWR VPWR registers\[29\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17377_ _15848_ _15853_ _15612_ VGND VGND VPWR VPWR _15854_ sky130_fd_sc_hd__o21ba_1
XFILLER_174_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_911 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19116_ registers\[36\]\[21\] registers\[37\]\[21\] registers\[38\]\[21\] registers\[39\]\[21\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__mux4_1
X_16328_ _14796_ _14833_ _14834_ _14799_ VGND VGND VPWR VPWR _14835_ sky130_fd_sc_hd__a22o_1
X_35162_ clknet_leaf_7_CLK _03276_ VGND VGND VPWR VPWR registers\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32374_ clknet_leaf_330_CLK _00488_ VGND VGND VPWR VPWR registers\[61\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34113_ clknet_leaf_259_CLK _02227_ VGND VGND VPWR VPWR registers\[35\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31325_ registers\[7\]\[23\] net16 _14157_ VGND VGND VPWR VPWR _14161_ sky130_fd_sc_hd__mux2_1
X_19047_ registers\[60\]\[19\] registers\[61\]\[19\] registers\[62\]\[19\] registers\[63\]\[19\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__mux4_1
X_16259_ registers\[12\]\[5\] registers\[13\]\[5\] registers\[14\]\[5\] registers\[15\]\[5\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14768_ sky130_fd_sc_hd__mux4_1
X_35093_ clknet_leaf_80_CLK _03207_ VGND VGND VPWR VPWR registers\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xoutput202 net202 VGND VGND VPWR VPWR D2[53] sky130_fd_sc_hd__buf_2
XFILLER_160_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput213 net213 VGND VGND VPWR VPWR D2[63] sky130_fd_sc_hd__buf_2
X_34044_ clknet_leaf_277_CLK _02158_ VGND VGND VPWR VPWR registers\[36\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31256_ _14124_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__clkbuf_1
Xoutput224 net224 VGND VGND VPWR VPWR D3[15] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR D3[25] sky130_fd_sc_hd__buf_2
XFILLER_47_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput246 net246 VGND VGND VPWR VPWR D3[35] sky130_fd_sc_hd__buf_2
XFILLER_47_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30207_ _13572_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__clkbuf_1
Xoutput257 net257 VGND VGND VPWR VPWR D3[45] sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR D3[55] sky130_fd_sc_hd__buf_2
XFILLER_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31187_ _14088_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__clkbuf_1
Xoutput279 net279 VGND VGND VPWR VPWR D3[7] sky130_fd_sc_hd__buf_2
XFILLER_86_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30138_ registers\[16\]\[37\] _13012_ _13528_ VGND VGND VPWR VPWR _13536_ sky130_fd_sc_hd__mux2_1
X_19949_ _06664_ _06667_ _06537_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__o21ba_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35995_ clknet_leaf_58_CLK _04109_ VGND VGND VPWR VPWR registers\[63\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22960_ net19 VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__clkbuf_4
X_34946_ clknet_leaf_205_CLK _03060_ VGND VGND VPWR VPWR registers\[22\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_30069_ registers\[16\]\[4\] _12943_ _13495_ VGND VGND VPWR VPWR _13500_ sky130_fd_sc_hd__mux2_1
XFILLER_110_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21911_ _08334_ _08573_ _08574_ _08338_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__a22o_1
XFILLER_228_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22891_ _09522_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34877_ clknet_leaf_186_CLK _02991_ VGND VGND VPWR VPWR registers\[23\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21842_ _08326_ _08506_ _08507_ _08332_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__a22o_1
X_24630_ _09561_ registers\[55\]\[22\] _10536_ VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__mux2_1
XFILLER_243_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33828_ clknet_leaf_471_CLK _01942_ VGND VGND VPWR VPWR registers\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_24561_ _09630_ registers\[56\]\[55\] _10495_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__mux2_1
X_21773_ registers\[48\]\[31\] registers\[49\]\[31\] registers\[50\]\[31\] registers\[51\]\[31\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__mux4_1
X_33759_ clknet_leaf_40_CLK _01873_ VGND VGND VPWR VPWR registers\[40\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26300_ _11453_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
X_20724_ registers\[4\]\[1\] registers\[5\]\[1\] registers\[6\]\[1\] registers\[7\]\[1\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__mux4_1
X_23512_ _09598_ registers\[19\]\[40\] _09914_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__mux2_1
X_27280_ _12000_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__clkbuf_1
X_24492_ _09561_ registers\[56\]\[22\] _10462_ VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__mux2_1
XFILLER_223_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23443_ _09878_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
X_26231_ _11417_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
X_20655_ _07343_ _07346_ _07351_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__a22o_1
X_35429_ clknet_leaf_461_CLK _03543_ VGND VGND VPWR VPWR registers\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_196_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26162_ _10747_ registers\[44\]\[8\] _11372_ VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__mux2_1
XFILLER_149_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23374_ registers\[39\]\[40\] _09775_ _09840_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__mux2_1
XFILLER_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20586_ _07284_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__buf_12
XFILLER_176_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22325_ registers\[44\]\[47\] registers\[45\]\[47\] registers\[46\]\[47\] registers\[47\]\[47\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__mux4_1
X_25113_ _10812_ registers\[52\]\[39\] _10794_ VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__mux2_1
XFILLER_165_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26093_ _11344_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
X_29921_ _13421_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__clkbuf_1
X_25044_ net9 VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__buf_2
X_22256_ registers\[36\]\[45\] registers\[37\]\[45\] registers\[38\]\[45\] registers\[39\]\[45\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__mux4_1
XFILLER_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21207_ _07287_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__buf_4
X_29852_ _13385_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_160_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_160_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_191_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22187_ registers\[32\]\[43\] registers\[33\]\[43\] registers\[34\]\[43\] registers\[35\]\[43\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__mux4_1
X_28803_ _11753_ registers\[25\]\[11\] _12801_ VGND VGND VPWR VPWR _12803_ sky130_fd_sc_hd__mux2_1
X_21138_ registers\[52\]\[13\] registers\[53\]\[13\] registers\[54\]\[13\] registers\[55\]\[13\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__mux4_1
X_29783_ registers\[1\]\[61\] _13062_ _13281_ VGND VGND VPWR VPWR _13349_ sky130_fd_sc_hd__mux2_1
X_26995_ _11846_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_1
X_28734_ _12766_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21069_ registers\[60\]\[11\] registers\[61\]\[11\] registers\[62\]\[11\] registers\[63\]\[11\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__mux4_1
X_25946_ _11267_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28665_ _12718_ VGND VGND VPWR VPWR _12730_ sky130_fd_sc_hd__buf_4
X_25877_ _11231_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27616_ _12178_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24828_ _09622_ registers\[54\]\[51\] _10642_ VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__mux2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28596_ _11816_ registers\[27\]\[41\] _12692_ VGND VGND VPWR VPWR _12694_ sky130_fd_sc_hd__mux2_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_12_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_12_0_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27547_ _11849_ registers\[35\]\[57\] _12133_ VGND VGND VPWR VPWR _12141_ sky130_fd_sc_hd__mux2_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24759_ _10607_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17300_ registers\[32\]\[35\] registers\[33\]\[35\] registers\[34\]\[35\] registers\[35\]\[35\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15779_ sky130_fd_sc_hd__mux4_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__buf_6
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27478_ _11780_ registers\[35\]\[24\] _12100_ VGND VGND VPWR VPWR _12105_ sky130_fd_sc_hd__mux2_1
XFILLER_203_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29217_ registers\[23\]\[53\] _13046_ _13040_ VGND VGND VPWR VPWR _13047_ sky130_fd_sc_hd__mux2_1
X_17231_ _15689_ _15696_ _15703_ _15712_ VGND VGND VPWR VPWR _15713_ sky130_fd_sc_hd__or4_4
X_26429_ _11521_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_27_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_27_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_196_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29148_ net25 VGND VGND VPWR VPWR _13000_ sky130_fd_sc_hd__clkbuf_4
X_17162_ _15637_ _15644_ _15645_ VGND VGND VPWR VPWR _15646_ sky130_fd_sc_hd__o21ba_1
XFILLER_196_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16113_ registers\[56\]\[1\] registers\[57\]\[1\] registers\[58\]\[1\] registers\[59\]\[1\]
+ _14530_ _14532_ VGND VGND VPWR VPWR _14626_ sky130_fd_sc_hd__mux4_1
X_29079_ net64 VGND VGND VPWR VPWR _12953_ sky130_fd_sc_hd__clkbuf_4
X_17093_ registers\[44\]\[29\] registers\[45\]\[29\] registers\[46\]\[29\] registers\[47\]\[29\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15578_ sky130_fd_sc_hd__mux4_1
XFILLER_196_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31110_ _14047_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16044_ _14490_ VGND VGND VPWR VPWR _14558_ sky130_fd_sc_hd__buf_4
XFILLER_143_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32090_ clknet_leaf_489_CLK _00003_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dfxtp_1
XFILLER_124_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31041_ _14011_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_151_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_151_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_151_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19803_ registers\[24\]\[40\] registers\[25\]\[40\] registers\[26\]\[40\] registers\[27\]\[40\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__mux4_1
XFILLER_170_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17995_ _14564_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__buf_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34800_ clknet_leaf_384_CLK _02914_ VGND VGND VPWR VPWR registers\[24\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_19734_ _06182_ _06457_ _06458_ _06185_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__a22o_1
X_16946_ registers\[40\]\[25\] registers\[41\]\[25\] registers\[42\]\[25\] registers\[43\]\[25\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15435_ sky130_fd_sc_hd__mux4_1
X_35780_ clknet_leaf_224_CLK _03894_ VGND VGND VPWR VPWR registers\[0\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_32992_ clknet_leaf_44_CLK _01106_ VGND VGND VPWR VPWR registers\[52\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31943_ _14485_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__clkbuf_1
X_19665_ _06187_ _06390_ _06391_ _06192_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__a22o_1
X_34731_ clknet_leaf_452_CLK _02845_ VGND VGND VPWR VPWR registers\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16877_ _15363_ _15368_ _15302_ VGND VGND VPWR VPWR _15369_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18616_ registers\[36\]\[7\] registers\[37\]\[7\] registers\[38\]\[7\] registers\[39\]\[7\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__mux4_1
XFILLER_77_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34662_ clknet_leaf_451_CLK _02776_ VGND VGND VPWR VPWR registers\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_19596_ _06321_ _06324_ _06194_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__o21ba_1
X_31874_ _14449_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33613_ clknet_leaf_76_CLK _01727_ VGND VGND VPWR VPWR registers\[43\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18547_ registers\[56\]\[5\] registers\[57\]\[5\] registers\[58\]\[5\] registers\[59\]\[5\]
+ _05272_ _05081_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux4_1
X_30825_ _09780_ registers\[11\]\[42\] _13895_ VGND VGND VPWR VPWR _13898_ sky130_fd_sc_hd__mux2_1
XFILLER_234_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34593_ clknet_leaf_8_CLK _02707_ VGND VGND VPWR VPWR registers\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33544_ clknet_leaf_251_CLK _01658_ VGND VGND VPWR VPWR registers\[44\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_18478_ registers\[36\]\[3\] registers\[37\]\[3\] registers\[38\]\[3\] registers\[39\]\[3\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__mux4_1
X_30756_ _13861_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17429_ registers\[4\]\[38\] registers\[5\]\[38\] registers\[6\]\[38\] registers\[7\]\[38\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _15905_ sky130_fd_sc_hd__mux4_1
X_33475_ clknet_leaf_255_CLK _01589_ VGND VGND VPWR VPWR registers\[45\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30687_ _13825_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35214_ clknet_leaf_112_CLK _03328_ VGND VGND VPWR VPWR registers\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_20440_ registers\[0\]\[59\] registers\[1\]\[59\] registers\[2\]\[59\] registers\[3\]\[59\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__mux4_1
XFILLER_14_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32426_ clknet_leaf_403_CLK _00540_ VGND VGND VPWR VPWR registers\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_36194_ clknet_leaf_98_CLK _00076_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35145_ clknet_leaf_218_CLK _03259_ VGND VGND VPWR VPWR registers\[1\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20371_ _07073_ _07076_ _06847_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__o21ba_1
XFILLER_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32357_ clknet_leaf_450_CLK _00471_ VGND VGND VPWR VPWR registers\[61\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_390_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_390_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22110_ _07329_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31308_ registers\[7\]\[15\] net7 _14146_ VGND VGND VPWR VPWR _14152_ sky130_fd_sc_hd__mux2_1
X_35076_ clknet_leaf_204_CLK _03190_ VGND VGND VPWR VPWR registers\[20\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_23090_ net12 VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__buf_4
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32288_ clknet_leaf_2_CLK _00402_ VGND VGND VPWR VPWR registers\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34027_ clknet_leaf_425_CLK _02141_ VGND VGND VPWR VPWR registers\[36\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_22041_ registers\[40\]\[39\] registers\[41\]\[39\] registers\[42\]\[39\] registers\[43\]\[39\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__mux4_1
XTAP_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_142_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_142_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31239_ _14115_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25800_ _11190_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
X_26780_ registers\[40\]\[44\] _10397_ _11702_ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__mux2_1
XFILLER_29_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35978_ clknet_leaf_158_CLK _04092_ VGND VGND VPWR VPWR registers\[6\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_23992_ _10170_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25731_ registers\[48\]\[61\] _10432_ _11085_ VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_11__f_CLK clknet_5_5_0_CLK VGND VGND VPWR VPWR clknet_6_11__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_34929_ clknet_leaf_385_CLK _03043_ VGND VGND VPWR VPWR registers\[22\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_22943_ _09556_ registers\[62\]\[20\] _09557_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28450_ _11805_ registers\[28\]\[36\] _12610_ VGND VGND VPWR VPWR _12617_ sky130_fd_sc_hd__mux2_1
X_25662_ registers\[48\]\[28\] _10363_ _11108_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__mux2_1
X_22874_ _09509_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27401_ _12064_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__clkbuf_1
X_24613_ _09544_ registers\[55\]\[14\] _10525_ VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__mux2_1
XFILLER_203_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28381_ _11736_ registers\[28\]\[3\] _12577_ VGND VGND VPWR VPWR _12581_ sky130_fd_sc_hd__mux2_1
X_21825_ _07361_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__buf_6
XFILLER_93_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25593_ registers\[4\]\[61\] _10432_ _11011_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__mux2_1
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27332_ registers\[36\]\[19\] _10344_ _12018_ VGND VGND VPWR VPWR _12028_ sky130_fd_sc_hd__mux2_1
X_24544_ _09613_ registers\[56\]\[47\] _10484_ VGND VGND VPWR VPWR _10492_ sky130_fd_sc_hd__mux2_1
X_21756_ _07315_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__buf_4
XFILLER_93_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20707_ registers\[44\]\[1\] registers\[45\]\[1\] registers\[46\]\[1\] registers\[47\]\[1\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__mux4_1
X_27263_ _11834_ registers\[37\]\[50\] _11991_ VGND VGND VPWR VPWR _11992_ sky130_fd_sc_hd__mux2_1
XFILLER_196_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21687_ _08357_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
X_24475_ _09544_ registers\[56\]\[14\] _10451_ VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__mux2_1
XFILLER_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29002_ _12907_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26214_ _11408_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
X_23426_ _09866_ _09868_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__nand2_8
XFILLER_196_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20638_ _07325_ _07330_ _07335_ _07336_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__a22o_1
XFILLER_32_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27194_ _11955_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26145_ _11371_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__buf_4
X_23357_ registers\[39\]\[32\] _09758_ _09829_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__mux2_1
X_20569_ registers\[28\]\[63\] registers\[29\]\[63\] registers\[30\]\[63\] registers\[31\]\[63\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__mux4_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_381_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_381_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22308_ _07366_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__buf_4
XFILLER_164_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23288_ _09787_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__clkbuf_1
X_26076_ _10796_ registers\[45\]\[31\] _11334_ VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29904_ registers\[18\]\[54\] _13048_ _13408_ VGND VGND VPWR VPWR _13413_ sky130_fd_sc_hd__mux2_1
X_22239_ _08615_ _08892_ _08893_ _08618_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__a22o_1
X_25027_ _10754_ registers\[52\]\[11\] _10752_ VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_133_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1705 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1716 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29835_ registers\[18\]\[21\] _12979_ _13375_ VGND VGND VPWR VPWR _13377_ sky130_fd_sc_hd__mux2_1
XTAP_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1727 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1738 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1749 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16800_ _15290_ _15291_ _15292_ _15293_ VGND VGND VPWR VPWR _15294_ sky130_fd_sc_hd__a22o_1
X_29766_ _13340_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__clkbuf_1
XTAP_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17780_ _14576_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__buf_6
XTAP_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26978_ _11729_ VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__buf_4
XFILLER_232_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16731_ _14952_ _15225_ _15226_ _14957_ VGND VGND VPWR VPWR _15227_ sky130_fd_sc_hd__a22o_1
X_28717_ _12757_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__clkbuf_1
X_25929_ _11258_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29697_ _13281_ VGND VGND VPWR VPWR _13304_ sky130_fd_sc_hd__buf_4
XFILLER_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19450_ registers\[24\]\[30\] registers\[25\]\[30\] registers\[26\]\[30\] registers\[27\]\[30\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__mux4_1
X_28648_ _12721_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__clkbuf_1
X_16662_ _15159_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18401_ _05148_ _05161_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o21ba_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19381_ _05839_ _06114_ _06115_ _05842_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__a22o_1
X_28579_ _11799_ registers\[27\]\[33\] _12681_ VGND VGND VPWR VPWR _12685_ sky130_fd_sc_hd__mux2_1
X_16593_ registers\[40\]\[15\] registers\[41\]\[15\] registers\[42\]\[15\] registers\[43\]\[15\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15092_ sky130_fd_sc_hd__mux4_1
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30610_ registers\[12\]\[4\] _12943_ _13780_ VGND VGND VPWR VPWR _13785_ sky130_fd_sc_hd__mux2_1
X_18332_ _05041_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__buf_12
XFILLER_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31590_ _14300_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ registers\[4\]\[63\] registers\[5\]\[63\] registers\[6\]\[63\] registers\[7\]\[63\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux4_1
XFILLER_124_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30541_ _13748_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17214_ _15692_ _15695_ _15620_ _15621_ VGND VGND VPWR VPWR _15696_ sky130_fd_sc_hd__o211a_1
X_33260_ clknet_leaf_365_CLK _01374_ VGND VGND VPWR VPWR registers\[48\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_30472_ _13712_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__clkbuf_1
X_18194_ _14587_ _04958_ _04959_ _14597_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__a22o_1
XFILLER_200_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32211_ clknet_leaf_332_CLK _00325_ VGND VGND VPWR VPWR registers\[9\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17145_ registers\[4\]\[30\] registers\[5\]\[30\] registers\[6\]\[30\] registers\[7\]\[30\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15629_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_372_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_372_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33191_ clknet_leaf_459_CLK _01305_ VGND VGND VPWR VPWR registers\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32142_ clknet_leaf_133_CLK _00256_ VGND VGND VPWR VPWR registers\[39\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_17076_ registers\[4\]\[28\] registers\[5\]\[28\] registers\[6\]\[28\] registers\[7\]\[28\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15562_ sky130_fd_sc_hd__mux4_1
XFILLER_226_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16027_ _14492_ VGND VGND VPWR VPWR _14541_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_124_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_124_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32073_ clknet_leaf_162_CLK _00251_ VGND VGND VPWR VPWR registers\[62\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35901_ clknet_leaf_305_CLK _04015_ VGND VGND VPWR VPWR registers\[7\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31024_ _14002_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35832_ clknet_leaf_332_CLK _03946_ VGND VGND VPWR VPWR registers\[8\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17978_ _14529_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__buf_6
XFILLER_242_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16929_ registers\[0\]\[24\] registers\[1\]\[24\] registers\[2\]\[24\] registers\[3\]\[24\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15419_ sky130_fd_sc_hd__mux4_1
X_19717_ _05092_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__clkbuf_4
X_32975_ clknet_leaf_172_CLK _01089_ VGND VGND VPWR VPWR registers\[52\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_35763_ clknet_leaf_383_CLK _03877_ VGND VGND VPWR VPWR registers\[0\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34714_ clknet_leaf_18_CLK _02828_ VGND VGND VPWR VPWR registers\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_31926_ _09802_ registers\[49\]\[52\] _14474_ VGND VGND VPWR VPWR _14477_ sky130_fd_sc_hd__mux2_1
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19648_ registers\[8\]\[36\] registers\[9\]\[36\] registers\[10\]\[36\] registers\[11\]\[36\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__mux4_1
XFILLER_246_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35694_ clknet_leaf_391_CLK _03808_ VGND VGND VPWR VPWR registers\[10\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34645_ clknet_leaf_95_CLK _02759_ VGND VGND VPWR VPWR registers\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_19579_ _06098_ _06306_ _06307_ _06102_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__a22o_1
XFILLER_59_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31857_ _14440_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21610_ registers\[28\]\[26\] registers\[29\]\[26\] registers\[30\]\[26\] registers\[31\]\[26\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__mux4_1
X_30808_ _09762_ registers\[11\]\[34\] _13884_ VGND VGND VPWR VPWR _13889_ sky130_fd_sc_hd__mux2_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22590_ registers\[12\]\[54\] registers\[13\]\[54\] registers\[14\]\[54\] registers\[15\]\[54\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__mux4_1
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34576_ clknet_leaf_118_CLK _02690_ VGND VGND VPWR VPWR registers\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_31788_ _14404_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_894 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21541_ registers\[20\]\[24\] registers\[21\]\[24\] registers\[22\]\[24\] registers\[23\]\[24\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__mux4_1
X_30739_ _09660_ registers\[11\]\[1\] _13851_ VGND VGND VPWR VPWR _13853_ sky130_fd_sc_hd__mux2_1
XFILLER_179_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33527_ clknet_leaf_340_CLK _01641_ VGND VGND VPWR VPWR registers\[44\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24260_ _10314_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21472_ _07377_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__buf_6
X_33458_ clknet_leaf_364_CLK _01572_ VGND VGND VPWR VPWR registers\[45\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23211_ registers\[9\]\[21\] _09702_ _09735_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__mux2_1
XFILLER_53_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20423_ _07106_ _07113_ _07120_ _07127_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__or4_1
X_32409_ clknet_leaf_21_CLK _00523_ VGND VGND VPWR VPWR registers\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24191_ _10275_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
X_36177_ clknet_leaf_92_CLK _00097_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_363_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_363_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33389_ clknet_leaf_344_CLK _01503_ VGND VGND VPWR VPWR registers\[46\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23142_ net10 VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__buf_4
X_20354_ _05060_ _07059_ _07060_ _05066_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__a22o_1
X_35128_ clknet_leaf_315_CLK _03242_ VGND VGND VPWR VPWR registers\[1\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27950_ registers\[32\]\[55\] _10420_ _12348_ VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__mux2_1
X_23073_ _09645_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_115_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_115_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35059_ clknet_leaf_412_CLK _03173_ VGND VGND VPWR VPWR registers\[20\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_20285_ _06784_ _06992_ _06993_ _06788_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__a22o_1
XTAP_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26901_ _11782_ registers\[3\]\[25\] _11772_ VGND VGND VPWR VPWR _11783_ sky130_fd_sc_hd__mux2_1
XFILLER_1_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22024_ registers\[0\]\[38\] registers\[1\]\[38\] registers\[2\]\[38\] registers\[3\]\[38\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__mux4_1
XFILLER_66_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27881_ registers\[32\]\[22\] _10351_ _12315_ VGND VGND VPWR VPWR _12318_ sky130_fd_sc_hd__mux2_1
XFILLER_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29620_ _13263_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__clkbuf_1
XTAP_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26832_ net34 VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29551_ _13227_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__clkbuf_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26763_ registers\[40\]\[36\] _10380_ _11691_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__mux2_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23975_ _09510_ registers\[5\]\[0\] _10161_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__mux2_1
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28502_ _11857_ registers\[28\]\[61\] _12576_ VGND VGND VPWR VPWR _12644_ sky130_fd_sc_hd__mux2_1
XFILLER_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25714_ _11144_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
X_29482_ _09788_ registers\[21\]\[46\] _13184_ VGND VGND VPWR VPWR _13191_ sky130_fd_sc_hd__mux2_1
X_22926_ net7 VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__buf_6
XFILLER_5_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26694_ registers\[40\]\[3\] _10311_ _11658_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__mux2_1
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28433_ _11788_ registers\[28\]\[28\] _12599_ VGND VGND VPWR VPWR _12608_ sky130_fd_sc_hd__mux2_1
XFILLER_231_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25645_ _11085_ VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__buf_4
X_22857_ _07385_ _09491_ _09492_ _07395_ VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__a22o_1
XFILLER_186_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28364_ _12571_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__clkbuf_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21808_ registers\[56\]\[32\] registers\[57\]\[32\] registers\[58\]\[32\] registers\[59\]\[32\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__mux4_1
X_25576_ _11070_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22788_ registers\[44\]\[61\] registers\[45\]\[61\] registers\[46\]\[61\] registers\[47\]\[61\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__mux4_1
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27315_ _12019_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__clkbuf_1
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24527_ _09596_ registers\[56\]\[39\] _10473_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__mux2_1
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28295_ _12535_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__clkbuf_1
X_21739_ registers\[8\]\[30\] registers\[9\]\[30\] registers\[10\]\[30\] registers\[11\]\[30\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__mux4_1
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27246_ _11818_ registers\[37\]\[42\] _11980_ VGND VGND VPWR VPWR _11983_ sky130_fd_sc_hd__mux2_1
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24458_ _09527_ registers\[56\]\[6\] _10440_ VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__mux2_1
XFILLER_8_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23409_ registers\[39\]\[57\] _09813_ _09851_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27177_ _11946_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_354_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_354_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24389_ registers\[57\]\[46\] _10401_ _10389_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__mux2_1
XFILLER_126_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26128_ _10848_ registers\[45\]\[56\] _11356_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_106_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_106_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26059_ _10779_ registers\[45\]\[23\] _11323_ VGND VGND VPWR VPWR _11327_ sky130_fd_sc_hd__mux2_1
X_18950_ _05693_ _05694_ _05695_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__a22o_1
XFILLER_4_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1502 _07349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17901_ _14527_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__buf_6
XFILLER_117_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18881_ _05626_ _05629_ _05494_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1513 _07974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1524 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1535 _09632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1546 _10426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ registers\[36\]\[50\] registers\[37\]\[50\] registers\[38\]\[50\] registers\[39\]\[50\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__mux4_1
XFILLER_239_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1557 _11513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29818_ registers\[18\]\[13\] _12962_ _13364_ VGND VGND VPWR VPWR _13368_ sky130_fd_sc_hd__mux2_1
XTAP_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1568 _12434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1579 _13921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17763_ registers\[56\]\[48\] registers\[57\]\[48\] registers\[58\]\[48\] registers\[59\]\[48\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__mux4_1
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29749_ _13331_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16714_ _14516_ VGND VGND VPWR VPWR _15210_ sky130_fd_sc_hd__clkbuf_4
X_19502_ _05088_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32760_ clknet_leaf_333_CLK _00874_ VGND VGND VPWR VPWR registers\[56\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17694_ registers\[60\]\[46\] registers\[61\]\[46\] registers\[62\]\[46\] registers\[63\]\[46\]
+ _04412_ _15893_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__mux4_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19433_ registers\[60\]\[30\] registers\[61\]\[30\] registers\[62\]\[30\] registers\[63\]\[30\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__mux4_1
X_31711_ registers\[59\]\[14\] net6 _14359_ VGND VGND VPWR VPWR _14364_ sky130_fd_sc_hd__mux2_1
X_16645_ _15139_ _15140_ _15141_ _15142_ VGND VGND VPWR VPWR _15143_ sky130_fd_sc_hd__a22o_1
X_32691_ clknet_leaf_363_CLK _00805_ VGND VGND VPWR VPWR registers\[57\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_34430_ clknet_leaf_182_CLK _02544_ VGND VGND VPWR VPWR registers\[30\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31642_ _14327_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19364_ _05092_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__clkbuf_8
X_16576_ registers\[0\]\[14\] registers\[1\]\[14\] registers\[2\]\[14\] registers\[3\]\[14\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15076_ sky130_fd_sc_hd__mux4_1
XFILLER_90_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18315_ _05041_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__buf_12
XFILLER_187_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34361_ clknet_leaf_60_CLK _02475_ VGND VGND VPWR VPWR registers\[31\]\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31573_ _14291_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19295_ registers\[8\]\[26\] registers\[9\]\[26\] registers\[10\]\[26\] registers\[11\]\[26\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__mux4_1
XFILLER_176_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36100_ clknet_leaf_236_CLK _04214_ VGND VGND VPWR VPWR registers\[59\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_33312_ clknet_leaf_31_CLK _01426_ VGND VGND VPWR VPWR registers\[47\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18246_ registers\[32\]\[63\] registers\[33\]\[63\] registers\[34\]\[63\] registers\[35\]\[63\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__mux4_1
XFILLER_176_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30524_ _13739_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34292_ clknet_leaf_349_CLK _02406_ VGND VGND VPWR VPWR registers\[32\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36031_ clknet_leaf_293_CLK _04145_ VGND VGND VPWR VPWR registers\[63\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_33243_ clknet_leaf_35_CLK _01357_ VGND VGND VPWR VPWR registers\[48\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_18177_ registers\[16\]\[60\] registers\[17\]\[60\] registers\[18\]\[60\] registers\[19\]\[60\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__mux4_1
X_30455_ _09817_ registers\[14\]\[59\] _13693_ VGND VGND VPWR VPWR _13703_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_345_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_345_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17128_ _14524_ VGND VGND VPWR VPWR _15612_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33174_ clknet_leaf_69_CLK _01288_ VGND VGND VPWR VPWR registers\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30386_ _09744_ registers\[14\]\[26\] _13660_ VGND VGND VPWR VPWR _13667_ sky130_fd_sc_hd__mux2_1
XFILLER_116_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32125_ clknet_leaf_393_CLK _00041_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dfxtp_1
X_17059_ _14543_ VGND VGND VPWR VPWR _15545_ sky130_fd_sc_hd__buf_4
XFILLER_104_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20070_ _05092_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__buf_4
X_32056_ clknet_leaf_332_CLK _00234_ VGND VGND VPWR VPWR registers\[62\]\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31007_ registers\[0\]\[0\] _12931_ _13993_ VGND VGND VPWR VPWR _13994_ sky130_fd_sc_hd__mux2_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35815_ clknet_leaf_460_CLK _03929_ VGND VGND VPWR VPWR registers\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20972_ _07657_ _07662_ _07370_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35746_ clknet_leaf_465_CLK _03860_ VGND VGND VPWR VPWR registers\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_23760_ _10047_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32958_ clknet_leaf_290_CLK _01072_ VGND VGND VPWR VPWR registers\[53\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22711_ _07276_ _09350_ _09351_ _07286_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__a22o_1
XFILLER_54_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31909_ _09784_ registers\[49\]\[44\] _14463_ VGND VGND VPWR VPWR _14468_ sky130_fd_sc_hd__mux2_1
X_23691_ _10009_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__clkbuf_1
X_35677_ clknet_leaf_484_CLK _03791_ VGND VGND VPWR VPWR registers\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_213_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32889_ clknet_leaf_287_CLK _01003_ VGND VGND VPWR VPWR registers\[54\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_25430_ _10991_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34628_ clknet_leaf_219_CLK _02742_ VGND VGND VPWR VPWR registers\[27\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_22642_ registers\[56\]\[56\] registers\[57\]\[56\] registers\[58\]\[56\] registers\[59\]\[56\]
+ _09223_ _09013_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__mux4_1
XFILLER_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22573_ _09148_ _09216_ _09217_ _09153_ VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__a22o_1
XFILLER_222_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25361_ _10955_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34559_ clknet_leaf_306_CLK _02673_ VGND VGND VPWR VPWR registers\[28\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27100_ _11807_ registers\[38\]\[37\] _11898_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__mux2_1
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24312_ registers\[57\]\[21\] _10349_ _10347_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__mux2_1
X_28080_ _12422_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21524_ registers\[60\]\[24\] registers\[61\]\[24\] registers\[62\]\[24\] registers\[63\]\[24\]
+ _08198_ _07992_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__mux4_1
X_25292_ _10918_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27031_ _11738_ registers\[38\]\[4\] _11865_ VGND VGND VPWR VPWR _11870_ sky130_fd_sc_hd__mux2_1
X_36229_ clknet_leaf_121_CLK _00114_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dfxtp_1
X_24243_ _10302_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21455_ registers\[56\]\[22\] registers\[57\]\[22\] registers\[58\]\[22\] registers\[59\]\[22\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_336_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_336_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20406_ registers\[52\]\[58\] registers\[53\]\[58\] registers\[54\]\[58\] registers\[55\]\[58\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__mux4_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24174_ _09577_ registers\[58\]\[30\] _10266_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__mux2_1
X_21386_ registers\[8\]\[20\] registers\[9\]\[20\] registers\[10\]\[20\] registers\[11\]\[20\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__mux4_1
XFILLER_190_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20337_ _06912_ _07042_ _07043_ _06917_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__a22o_1
XFILLER_135_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23125_ registers\[39\]\[12\] _09683_ _09679_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__mux2_1
X_28982_ registers\[24\]\[32\] _10372_ _12894_ VGND VGND VPWR VPWR _12897_ sky130_fd_sc_hd__mux2_1
XFILLER_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23056_ net53 VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__buf_6
X_27933_ registers\[32\]\[47\] _10403_ _12337_ VGND VGND VPWR VPWR _12345_ sky130_fd_sc_hd__mux2_1
X_20268_ _06974_ _06977_ _06880_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__o21ba_1
XTAP_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22007_ _08664_ _08667_ _08397_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__o21ba_1
XTAP_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27864_ registers\[32\]\[14\] _10334_ _12304_ VGND VGND VPWR VPWR _12309_ sky130_fd_sc_hd__mux2_1
X_20199_ _06889_ _06896_ _06903_ _06910_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__or4_2
XFILLER_163_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26815_ registers\[40\]\[61\] _10432_ _11657_ VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__mux2_1
XTAP_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29603_ _13254_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27795_ _12272_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__clkbuf_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29534_ _13218_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__clkbuf_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26746_ registers\[40\]\[28\] _10363_ _11680_ VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23958_ _09634_ registers\[60\]\[57\] _10144_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__mux2_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_900 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_911 _09708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_922 _09791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22909_ _09534_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29465_ _09771_ registers\[21\]\[38\] _13173_ VGND VGND VPWR VPWR _13182_ sky130_fd_sc_hd__mux2_1
X_26677_ _10856_ registers\[41\]\[60\] _11585_ VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__mux2_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_933 _10016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_944 _10344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23889_ _09565_ registers\[60\]\[24\] _10111_ VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__mux2_1
X_28416_ _12576_ VGND VGND VPWR VPWR _12599_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_955 _10586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16430_ _14553_ VGND VGND VPWR VPWR _14934_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25628_ _11099_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_966 _10864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_977 _11229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29396_ _09668_ registers\[21\]\[5\] _13140_ VGND VGND VPWR VPWR _13146_ sky130_fd_sc_hd__mux2_1
XFILLER_108_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_988 _11729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_999 _11820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28347_ registers\[2\]\[51\] _10412_ _12561_ VGND VGND VPWR VPWR _12563_ sky130_fd_sc_hd__mux2_1
XFILLER_188_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16361_ _14516_ VGND VGND VPWR VPWR _14867_ sky130_fd_sc_hd__clkbuf_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25559_ _11061_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18100_ _04683_ _04867_ _04868_ _04686_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a22o_1
XFILLER_212_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19080_ registers\[60\]\[20\] registers\[61\]\[20\] registers\[62\]\[20\] registers\[63\]\[20\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__mux4_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _14796_ _14797_ _14798_ _14799_ VGND VGND VPWR VPWR _14800_ sky130_fd_sc_hd__a22o_1
X_28278_ _12526_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__clkbuf_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18031_ _04637_ _04801_ _04802_ _04642_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a22o_1
XFILLER_205_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27229_ _11801_ registers\[37\]\[34\] _11969_ VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__mux2_1
XFILLER_185_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_327_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_327_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30240_ registers\[15\]\[21\] _12979_ _13588_ VGND VGND VPWR VPWR _13590_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30171_ _13553_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19982_ _06676_ _06683_ _06692_ _06699_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__or4_4
XFILLER_207_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18933_ registers\[48\]\[16\] registers\[49\]\[16\] registers\[50\]\[16\] registers\[51\]\[16\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__mux4_1
XANTENNA_1310 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1321 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1332 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33930_ clknet_leaf_158_CLK _02044_ VGND VGND VPWR VPWR registers\[38\]\[60\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1343 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18864_ _05547_ _05611_ _05612_ _05550_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__a22o_1
XANTENNA_1354 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1365 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1376 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17815_ _04486_ _04591_ _04592_ _04489_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__a22o_1
XANTENNA_1387 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33861_ clknet_leaf_224_CLK _01975_ VGND VGND VPWR VPWR registers\[3\]\[55\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1398 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18795_ _05540_ _05543_ _05544_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__a22o_1
XTAP_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35600_ clknet_leaf_135_CLK _03714_ VGND VGND VPWR VPWR registers\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17746_ registers\[16\]\[47\] registers\[17\]\[47\] registers\[18\]\[47\] registers\[19\]\[47\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__mux4_1
X_32812_ clknet_leaf_373_CLK _00926_ VGND VGND VPWR VPWR registers\[55\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33792_ clknet_leaf_272_CLK _01906_ VGND VGND VPWR VPWR registers\[40\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35531_ clknet_leaf_150_CLK _03645_ VGND VGND VPWR VPWR registers\[13\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_17677_ _04289_ _04457_ _04458_ _04292_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__a22o_1
X_32743_ clknet_leaf_436_CLK _00857_ VGND VGND VPWR VPWR registers\[56\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19416_ _05844_ _06148_ _06149_ _05849_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__a22o_1
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16628_ registers\[44\]\[16\] registers\[45\]\[16\] registers\[46\]\[16\] registers\[47\]\[16\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15126_ sky130_fd_sc_hd__mux4_1
X_35462_ clknet_leaf_211_CLK _03576_ VGND VGND VPWR VPWR registers\[14\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_32674_ clknet_leaf_441_CLK _00788_ VGND VGND VPWR VPWR registers\[57\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34413_ clknet_leaf_403_CLK _02527_ VGND VGND VPWR VPWR registers\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_31625_ _14318_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__clkbuf_1
X_19347_ _06082_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_1
X_16559_ registers\[40\]\[14\] registers\[41\]\[14\] registers\[42\]\[14\] registers\[43\]\[14\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15059_ sky130_fd_sc_hd__mux4_1
X_35393_ clknet_leaf_238_CLK _03507_ VGND VGND VPWR VPWR registers\[15\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31556_ _14282_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__clkbuf_1
X_34344_ clknet_leaf_454_CLK _02458_ VGND VGND VPWR VPWR registers\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_19278_ registers\[40\]\[26\] registers\[41\]\[26\] registers\[42\]\[26\] registers\[43\]\[26\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__mux4_1
XFILLER_104_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18229_ registers\[8\]\[62\] registers\[9\]\[62\] registers\[10\]\[62\] registers\[11\]\[62\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__mux4_1
X_30507_ _13730_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34275_ clknet_leaf_56_CLK _02389_ VGND VGND VPWR VPWR registers\[32\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_318_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_318_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31487_ _09766_ registers\[6\]\[36\] _14239_ VGND VGND VPWR VPWR _14246_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33226_ clknet_leaf_156_CLK _01340_ VGND VGND VPWR VPWR registers\[4\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_36014_ clknet_leaf_370_CLK _04128_ VGND VGND VPWR VPWR registers\[63\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_21240_ _07917_ _07922_ _07719_ _07720_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__o211a_1
X_30438_ _13694_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33157_ clknet_leaf_259_CLK _01271_ VGND VGND VPWR VPWR registers\[50\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_21171_ registers\[60\]\[14\] registers\[61\]\[14\] registers\[62\]\[14\] registers\[63\]\[14\]
+ _07855_ _07649_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30369_ _09695_ registers\[14\]\[18\] _13649_ VGND VGND VPWR VPWR _13658_ sky130_fd_sc_hd__mux2_1
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20122_ _06530_ _06834_ _06835_ _06535_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__a22o_1
X_32108_ clknet_leaf_483_CLK _00023_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dfxtp_1
X_33088_ clknet_leaf_269_CLK _01202_ VGND VGND VPWR VPWR registers\[51\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24930_ _10697_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
X_20053_ _06768_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
X_32039_ clknet_leaf_437_CLK _00217_ VGND VGND VPWR VPWR registers\[62\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24861_ _10661_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26600_ _10779_ registers\[41\]\[23\] _11608_ VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__mux2_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23812_ _09624_ registers\[29\]\[52\] _10072_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__mux2_1
XFILLER_85_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27580_ _12159_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24792_ _09586_ registers\[54\]\[34\] _10620_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__mux2_1
XFILLER_2_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_207 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26531_ _10846_ registers\[42\]\[55\] _11569_ VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__mux2_1
XFILLER_213_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_218 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35729_ clknet_leaf_109_CLK _03843_ VGND VGND VPWR VPWR registers\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_23743_ _10038_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20955_ _07285_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__clkbuf_4
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29250_ _13068_ VGND VGND VPWR VPWR _13069_ sky130_fd_sc_hd__buf_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26462_ _10777_ registers\[42\]\[22\] _11536_ VGND VGND VPWR VPWR _11539_ sky130_fd_sc_hd__mux2_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23674_ registers\[61\]\[52\] _09802_ _09998_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__mux2_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20886_ _07325_ _07575_ _07578_ _07336_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__a22o_1
XFILLER_41_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28201_ _11826_ registers\[30\]\[46\] _12479_ VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__mux2_1
XFILLER_13_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25413_ _10817_ registers\[50\]\[41\] _10981_ VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__mux2_1
X_22625_ _09265_ _09268_ _09102_ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__o21ba_1
X_29181_ _13022_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26393_ _11502_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__clkbuf_1
X_28132_ _11757_ registers\[30\]\[13\] _12446_ VGND VGND VPWR VPWR _12450_ sky130_fd_sc_hd__mux2_1
XFILLER_167_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25344_ _10946_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__clkbuf_1
X_22556_ _07303_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__buf_6
XFILLER_22_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28063_ _12413_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_1
X_21507_ registers\[20\]\[23\] registers\[21\]\[23\] registers\[22\]\[23\] registers\[23\]\[23\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_309_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_309_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25275_ _10814_ registers\[51\]\[40\] _10909_ VGND VGND VPWR VPWR _10910_ sky130_fd_sc_hd__mux2_1
X_22487_ _08953_ _09133_ _09134_ _08956_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__a22o_1
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27014_ net59 VGND VGND VPWR VPWR _11859_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24226_ _09630_ registers\[58\]\[55\] _10288_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__mux2_1
XFILLER_170_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21438_ _08080_ _08114_ _08115_ _08085_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__a22o_1
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24157_ _09561_ registers\[58\]\[22\] _10255_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__mux2_1
X_21369_ _07776_ _08046_ _08047_ _07781_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__a22o_1
XFILLER_107_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23108_ net62 VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__buf_4
XFILLER_1_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24088_ _09628_ registers\[5\]\[54\] _10216_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__mux2_1
XFILLER_174_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28965_ registers\[24\]\[24\] _10355_ _12883_ VGND VGND VPWR VPWR _12888_ sky130_fd_sc_hd__mux2_1
XFILLER_231_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23039_ _09622_ registers\[62\]\[51\] _09620_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__mux2_1
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27916_ registers\[32\]\[39\] _10386_ _12326_ VGND VGND VPWR VPWR _12336_ sky130_fd_sc_hd__mux2_1
X_28896_ _12851_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__clkbuf_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27847_ registers\[32\]\[6\] _10317_ _12293_ VGND VGND VPWR VPWR _12300_ sky130_fd_sc_hd__mux2_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ registers\[8\]\[43\] registers\[9\]\[43\] registers\[10\]\[43\] registers\[11\]\[43\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__mux4_1
XFILLER_218_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ registers\[48\]\[6\] registers\[49\]\[6\] registers\[50\]\[6\] registers\[51\]\[6\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux4_1
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27778_ _12263_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__clkbuf_1
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _04313_ _04316_ _15963_ _15964_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__o211a_1
X_29517_ _09825_ registers\[21\]\[63\] _13139_ VGND VGND VPWR VPWR _13209_ sky130_fd_sc_hd__mux2_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26729_ _11657_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__buf_4
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_730 _07352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_741 _07363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_752 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29448_ _13139_ VGND VGND VPWR VPWR _13173_ sky130_fd_sc_hd__buf_4
X_17462_ _15830_ _15935_ _15936_ _15833_ VGND VGND VPWR VPWR _15937_ sky130_fd_sc_hd__a22o_1
XFILLER_229_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_763 _07571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_774 _08089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19201_ _05693_ _05939_ _05940_ _05696_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__a22o_1
X_16413_ _14917_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_785 _08775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_796 _08905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29379_ _13136_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17393_ registers\[16\]\[37\] registers\[17\]\[37\] registers\[18\]\[37\] registers\[19\]\[37\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _15870_ sky130_fd_sc_hd__mux4_1
XFILLER_186_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31410_ _10159_ _10585_ VGND VGND VPWR VPWR _14205_ sky130_fd_sc_hd__nand2_8
X_19132_ _05870_ _05873_ _05837_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__o21ba_1
X_16344_ _14648_ _14848_ _14849_ _14653_ VGND VGND VPWR VPWR _14850_ sky130_fd_sc_hd__a22o_1
XFILLER_185_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32390_ clknet_leaf_198_CLK _00504_ VGND VGND VPWR VPWR registers\[61\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19063_ _05501_ _05805_ _05806_ _05506_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__a22o_1
X_31341_ _14169_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__clkbuf_1
X_16275_ registers\[44\]\[6\] registers\[45\]\[6\] registers\[46\]\[6\] registers\[47\]\[6\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14783_ sky130_fd_sc_hd__mux4_1
XFILLER_158_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1030 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18014_ _04540_ _04784_ _04785_ _04546_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a22o_1
XFILLER_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34060_ clknet_leaf_172_CLK _02174_ VGND VGND VPWR VPWR registers\[36\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_31272_ _14132_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33011_ clknet_leaf_360_CLK _01125_ VGND VGND VPWR VPWR registers\[52\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_30223_ registers\[15\]\[13\] _12962_ _13577_ VGND VGND VPWR VPWR _13581_ sky130_fd_sc_hd__mux2_1
XFILLER_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30154_ _13544_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19965_ _06679_ _06682_ _06512_ _06513_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__o211a_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18916_ registers\[24\]\[15\] registers\[25\]\[15\] registers\[26\]\[15\] registers\[27\]\[15\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__mux4_1
XTAP_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34962_ clknet_leaf_100_CLK _03076_ VGND VGND VPWR VPWR registers\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_30085_ _13508_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1140 _14632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19896_ registers\[60\]\[43\] registers\[61\]\[43\] registers\[62\]\[43\] registers\[63\]\[43\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__mux4_1
XANTENNA_1151 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1162 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33913_ clknet_leaf_281_CLK _02027_ VGND VGND VPWR VPWR registers\[38\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1173 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18847_ registers\[4\]\[13\] registers\[5\]\[13\] registers\[6\]\[13\] registers\[7\]\[13\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__mux4_1
X_34893_ clknet_leaf_145_CLK _03007_ VGND VGND VPWR VPWR registers\[23\]\[63\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1184 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1195 _15915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33844_ clknet_leaf_415_CLK _01958_ VGND VGND VPWR VPWR registers\[3\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_18778_ _05350_ _05528_ _05529_ _05353_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__a22o_1
XFILLER_247_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17729_ _04340_ _04505_ _04508_ _04343_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a22o_1
XFILLER_247_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30987_ registers\[10\]\[55\] _13050_ _13977_ VGND VGND VPWR VPWR _13983_ sky130_fd_sc_hd__mux2_1
X_33775_ clknet_leaf_347_CLK _01889_ VGND VGND VPWR VPWR registers\[40\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35514_ clknet_leaf_303_CLK _03628_ VGND VGND VPWR VPWR registers\[13\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20740_ registers\[32\]\[2\] registers\[33\]\[2\] registers\[34\]\[2\] registers\[35\]\[2\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__mux4_1
XFILLER_208_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32726_ clknet_leaf_65_CLK _00840_ VGND VGND VPWR VPWR registers\[56\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20671_ _07369_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__buf_2
X_35445_ clknet_leaf_323_CLK _03559_ VGND VGND VPWR VPWR registers\[14\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_32657_ clknet_leaf_74_CLK _00771_ VGND VGND VPWR VPWR registers\[57\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_95_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22410_ registers\[8\]\[49\] registers\[9\]\[49\] registers\[10\]\[49\] registers\[11\]\[49\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__mux4_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31608_ _14309_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__clkbuf_1
X_32588_ clknet_leaf_144_CLK _00702_ VGND VGND VPWR VPWR registers\[5\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_23390_ registers\[39\]\[48\] _09793_ _09840_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__mux2_1
X_35376_ clknet_leaf_375_CLK _03490_ VGND VGND VPWR VPWR registers\[15\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34327_ clknet_leaf_98_CLK _02441_ VGND VGND VPWR VPWR registers\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_22341_ registers\[12\]\[47\] registers\[13\]\[47\] registers\[14\]\[47\] registers\[15\]\[47\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__mux4_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31539_ _09821_ registers\[6\]\[61\] _14205_ VGND VGND VPWR VPWR _14273_ sky130_fd_sc_hd__mux2_1
XFILLER_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22272_ registers\[4\]\[45\] registers\[5\]\[45\] registers\[6\]\[45\] registers\[7\]\[45\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__mux4_1
X_25060_ net15 VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__buf_2
X_34258_ clknet_leaf_122_CLK _02372_ VGND VGND VPWR VPWR registers\[32\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24011_ _10180_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
X_21223_ _07883_ _07890_ _07899_ _07906_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__or4_2
X_33209_ clknet_leaf_315_CLK _01323_ VGND VGND VPWR VPWR registers\[4\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_34189_ clknet_leaf_170_CLK _02303_ VGND VGND VPWR VPWR registers\[34\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21154_ registers\[20\]\[13\] registers\[21\]\[13\] registers\[22\]\[13\] registers\[23\]\[13\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__mux4_1
XFILLER_104_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20105_ _06776_ _06817_ _06818_ _06782_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__a22o_1
XFILLER_144_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28750_ _11834_ registers\[26\]\[50\] _12774_ VGND VGND VPWR VPWR _12775_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21085_ _07737_ _07771_ _07772_ _07742_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__a22o_1
X_25962_ _10817_ registers\[46\]\[41\] _11274_ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27701_ _12223_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__clkbuf_1
X_20036_ _06441_ _06750_ _06751_ _06445_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__a22o_1
X_24913_ _10688_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28681_ _12738_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25893_ _11239_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27632_ registers\[34\]\[32\] _10372_ _12184_ VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__mux2_1
X_24844_ _09638_ registers\[54\]\[59\] _10642_ VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__mux2_1
XFILLER_73_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27563_ _09653_ _12149_ VGND VGND VPWR VPWR _12150_ sky130_fd_sc_hd__nor2_8
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24775_ _09569_ registers\[54\]\[26\] _10609_ VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__mux2_1
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21987_ _08610_ _08647_ _08648_ _08613_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__a22o_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29302_ _13096_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__clkbuf_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26514_ _10829_ registers\[42\]\[47\] _11558_ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__mux2_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _09538_ registers\[29\]\[11\] _10028_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__mux2_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _07386_ _07628_ _07629_ _07396_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__a22o_1
XFILLER_15_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27494_ _12113_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__clkbuf_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29233_ _13057_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__clkbuf_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26445_ _10760_ registers\[42\]\[14\] _11525_ VGND VGND VPWR VPWR _11530_ sky130_fd_sc_hd__mux2_1
X_23657_ registers\[61\]\[44\] _09784_ _09987_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__mux2_1
XFILLER_42_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _07559_ _07562_ _07399_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_86_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_86_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22608_ registers\[44\]\[55\] registers\[45\]\[55\] registers\[46\]\[55\] registers\[47\]\[55\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__mux4_1
XFILLER_161_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29164_ registers\[23\]\[36\] _13010_ _12998_ VGND VGND VPWR VPWR _13011_ sky130_fd_sc_hd__mux2_1
XFILLER_53_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26376_ _11493_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23588_ registers\[61\]\[11\] _09681_ _09954_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__mux2_1
XFILLER_169_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28115_ _11740_ registers\[30\]\[5\] _12435_ VGND VGND VPWR VPWR _12441_ sky130_fd_sc_hd__mux2_1
X_25327_ _10728_ registers\[50\]\[0\] _10937_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__mux2_1
XFILLER_168_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22539_ registers\[40\]\[53\] registers\[41\]\[53\] registers\[42\]\[53\] registers\[43\]\[53\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__mux4_1
X_29095_ net6 VGND VGND VPWR VPWR _12964_ sky130_fd_sc_hd__buf_4
XFILLER_167_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16060_ _14573_ VGND VGND VPWR VPWR _14574_ sky130_fd_sc_hd__buf_6
X_28046_ _12404_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_1
X_25258_ _10798_ registers\[51\]\[32\] _10898_ VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__mux2_1
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24209_ _09613_ registers\[58\]\[47\] _10277_ VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__mux2_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25189_ _09868_ _10512_ VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__nand2_8
XFILLER_155_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29997_ registers\[17\]\[34\] _13006_ _13457_ VGND VGND VPWR VPWR _13462_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19750_ registers\[56\]\[39\] registers\[57\]\[39\] registers\[58\]\[39\] registers\[59\]\[39\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__mux4_1
XFILLER_111_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16962_ registers\[8\]\[25\] registers\[9\]\[25\] registers\[10\]\[25\] registers\[11\]\[25\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15451_ sky130_fd_sc_hd__mux4_1
X_28948_ registers\[24\]\[16\] _10338_ _12872_ VGND VGND VPWR VPWR _12879_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_10_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_231_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18701_ registers\[12\]\[9\] registers\[13\]\[9\] registers\[14\]\[9\] registers\[15\]\[9\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19681_ registers\[60\]\[37\] registers\[61\]\[37\] registers\[62\]\[37\] registers\[63\]\[37\]
+ _06305_ _06099_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__mux4_1
X_16893_ _15380_ _15383_ _15277_ _15278_ VGND VGND VPWR VPWR _15384_ sky130_fd_sc_hd__o211a_1
XFILLER_103_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28879_ _12842_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18632_ _05384_ _05387_ _05134_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__o21ba_1
X_30910_ _13942_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__clkbuf_1
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31890_ _09764_ registers\[49\]\[35\] _14452_ VGND VGND VPWR VPWR _14458_ sky130_fd_sc_hd__mux2_1
XFILLER_209_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30841_ _13850_ VGND VGND VPWR VPWR _13906_ sky130_fd_sc_hd__buf_4
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18563_ registers\[24\]\[5\] registers\[25\]\[5\] registers\[26\]\[5\] registers\[27\]\[5\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__mux4_1
XFILLER_224_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17514_ _14613_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__buf_2
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18494_ registers\[4\]\[3\] registers\[5\]\[3\] registers\[6\]\[3\] registers\[7\]\[3\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__mux4_1
X_33560_ clknet_leaf_90_CLK _01674_ VGND VGND VPWR VPWR registers\[43\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_30772_ _09693_ registers\[11\]\[17\] _13862_ VGND VGND VPWR VPWR _13870_ sky130_fd_sc_hd__mux2_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_560 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_571 _04892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32511_ clknet_leaf_291_CLK _00625_ VGND VGND VPWR VPWR registers\[60\]\[49\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_582 _05053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _15677_ _15916_ _15919_ _15682_ VGND VGND VPWR VPWR _15920_ sky130_fd_sc_hd__a22o_1
X_33491_ clknet_leaf_129_CLK _01605_ VGND VGND VPWR VPWR registers\[44\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_593 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_77_CLK sky130_fd_sc_hd__clkbuf_16
X_32442_ clknet_leaf_184_CLK _00556_ VGND VGND VPWR VPWR registers\[29\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_35230_ clknet_leaf_3_CLK _03344_ VGND VGND VPWR VPWR registers\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17376_ _15684_ _15849_ _15852_ _15687_ VGND VGND VPWR VPWR _15853_ sky130_fd_sc_hd__a22o_1
XFILLER_14_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16327_ registers\[0\]\[7\] registers\[1\]\[7\] registers\[2\]\[7\] registers\[3\]\[7\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14834_ sky130_fd_sc_hd__mux4_1
XFILLER_140_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19115_ registers\[44\]\[21\] registers\[45\]\[21\] registers\[46\]\[21\] registers\[47\]\[21\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__mux4_2
XFILLER_174_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35161_ clknet_leaf_6_CLK _03275_ VGND VGND VPWR VPWR registers\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_32373_ clknet_leaf_353_CLK _00487_ VGND VGND VPWR VPWR registers\[61\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34112_ clknet_leaf_270_CLK _02226_ VGND VGND VPWR VPWR registers\[35\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_31324_ _14160_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__clkbuf_1
X_19046_ _05747_ _05788_ _05789_ _05753_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__a22o_1
X_16258_ _14558_ _14765_ _14766_ _14568_ VGND VGND VPWR VPWR _14767_ sky130_fd_sc_hd__a22o_1
X_35092_ clknet_leaf_80_CLK _03206_ VGND VGND VPWR VPWR registers\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput203 net203 VGND VGND VPWR VPWR D2[54] sky130_fd_sc_hd__buf_2
XFILLER_86_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31255_ registers\[8\]\[54\] net50 _14119_ VGND VGND VPWR VPWR _14124_ sky130_fd_sc_hd__mux2_1
X_34043_ clknet_leaf_282_CLK _02157_ VGND VGND VPWR VPWR registers\[36\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_16189_ registers\[0\]\[3\] registers\[1\]\[3\] registers\[2\]\[3\] registers\[3\]\[3\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14700_ sky130_fd_sc_hd__mux4_1
XFILLER_160_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 net214 VGND VGND VPWR VPWR D2[6] sky130_fd_sc_hd__buf_2
XFILLER_154_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput225 net225 VGND VGND VPWR VPWR D3[16] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR D3[26] sky130_fd_sc_hd__buf_2
X_30206_ registers\[15\]\[5\] _12945_ _13566_ VGND VGND VPWR VPWR _13572_ sky130_fd_sc_hd__mux2_1
Xoutput247 net247 VGND VGND VPWR VPWR D3[36] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR D3[46] sky130_fd_sc_hd__buf_2
XFILLER_142_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31186_ registers\[8\]\[21\] net14 _14086_ VGND VGND VPWR VPWR _14088_ sky130_fd_sc_hd__mux2_1
Xoutput269 net269 VGND VGND VPWR VPWR D3[56] sky130_fd_sc_hd__buf_2
XFILLER_173_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30137_ _13535_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__clkbuf_1
X_19948_ _06530_ _06665_ _06666_ _06535_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__a22o_1
X_35994_ clknet_leaf_62_CLK _04108_ VGND VGND VPWR VPWR registers\[63\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34945_ clknet_leaf_202_CLK _03059_ VGND VGND VPWR VPWR registers\[22\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30068_ _13499_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__clkbuf_1
X_19879_ _05127_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__buf_4
XFILLER_214_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21910_ registers\[52\]\[35\] registers\[53\]\[35\] registers\[54\]\[35\] registers\[55\]\[35\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__mux4_1
XFILLER_216_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22890_ _09521_ registers\[62\]\[3\] _09515_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__mux2_1
X_34876_ clknet_leaf_188_CLK _02990_ VGND VGND VPWR VPWR registers\[23\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33827_ clknet_leaf_471_CLK _01941_ VGND VGND VPWR VPWR registers\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_21841_ registers\[48\]\[33\] registers\[49\]\[33\] registers\[50\]\[33\] registers\[51\]\[33\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__mux4_1
XFILLER_3_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24560_ _10500_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
X_21772_ registers\[56\]\[31\] registers\[57\]\[31\] registers\[58\]\[31\] registers\[59\]\[31\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__mux4_1
X_33758_ clknet_leaf_27_CLK _01872_ VGND VGND VPWR VPWR registers\[40\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23511_ _09869_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__clkbuf_8
X_20723_ registers\[12\]\[1\] registers\[13\]\[1\] registers\[14\]\[1\] registers\[15\]\[1\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__mux4_1
X_32709_ clknet_leaf_264_CLK _00823_ VGND VGND VPWR VPWR registers\[57\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24491_ _10464_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_68_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_68_CLK sky130_fd_sc_hd__clkbuf_16
X_33689_ clknet_leaf_90_CLK _01803_ VGND VGND VPWR VPWR registers\[41\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_26230_ _10814_ registers\[44\]\[40\] _11416_ VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__mux2_1
XFILLER_168_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23442_ _09529_ registers\[19\]\[7\] _09870_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__mux2_1
X_35428_ clknet_leaf_467_CLK _03542_ VGND VGND VPWR VPWR registers\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20654_ _07352_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__buf_4
XFILLER_221_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26161_ _11380_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20585_ net73 net74 VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__nor2_4
X_23373_ _09657_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__buf_4
X_35359_ clknet_leaf_482_CLK _03473_ VGND VGND VPWR VPWR registers\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_25112_ net33 VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__buf_2
X_22324_ _08805_ _08974_ _08975_ _08810_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__a22o_1
XFILLER_137_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26092_ _10812_ registers\[45\]\[39\] _11334_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_34__f_CLK clknet_5_17_0_CLK VGND VGND VPWR VPWR clknet_6_34__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_29920_ registers\[18\]\[62\] _13064_ _13352_ VGND VGND VPWR VPWR _13421_ sky130_fd_sc_hd__mux2_1
XFILLER_124_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25043_ _10765_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
X_22255_ registers\[44\]\[45\] registers\[45\]\[45\] registers\[46\]\[45\] registers\[47\]\[45\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__mux4_1
XFILLER_219_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21206_ _07886_ _07889_ _07719_ _07720_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__o211a_1
XFILLER_195_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22186_ registers\[40\]\[43\] registers\[41\]\[43\] registers\[42\]\[43\] registers\[43\]\[43\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__mux4_1
X_29851_ registers\[18\]\[29\] _12995_ _13375_ VGND VGND VPWR VPWR _13385_ sky130_fd_sc_hd__mux2_1
XFILLER_152_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28802_ _12802_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21137_ registers\[60\]\[13\] registers\[61\]\[13\] registers\[62\]\[13\] registers\[63\]\[13\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__mux4_1
XFILLER_48_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29782_ _13348_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__clkbuf_1
X_26994_ _11845_ registers\[3\]\[55\] _11835_ VGND VGND VPWR VPWR _11846_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21068_ _07640_ _07754_ _07755_ _07646_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__a22o_1
X_25945_ _10800_ registers\[46\]\[33\] _11263_ VGND VGND VPWR VPWR _11267_ sky130_fd_sc_hd__mux2_1
X_28733_ _11818_ registers\[26\]\[42\] _12763_ VGND VGND VPWR VPWR _12766_ sky130_fd_sc_hd__mux2_1
XFILLER_171_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20019_ _06732_ _06735_ _06537_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__o21ba_1
X_28664_ _12729_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25876_ _10728_ registers\[46\]\[0\] _11230_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__mux2_1
XFILLER_171_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24827_ _10643_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27615_ registers\[34\]\[24\] _10355_ _12173_ VGND VGND VPWR VPWR _12178_ sky130_fd_sc_hd__mux2_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28595_ _12693_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__clkbuf_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27546_ _12140_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__clkbuf_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_802 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24758_ _09552_ registers\[54\]\[18\] _10598_ VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__mux2_1
XFILLER_76_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23709_ _09521_ registers\[29\]\[3\] _10017_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__mux2_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27477_ _12104_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24689_ _09619_ registers\[55\]\[50\] _10569_ VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_59_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _15706_ _15711_ _15645_ VGND VGND VPWR VPWR _15712_ sky130_fd_sc_hd__o21ba_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29216_ net49 VGND VGND VPWR VPWR _13046_ sky130_fd_sc_hd__buf_4
X_26428_ _10743_ registers\[42\]\[6\] _11514_ VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__mux2_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29147_ _12999_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__clkbuf_1
X_17161_ _14613_ VGND VGND VPWR VPWR _15645_ sky130_fd_sc_hd__buf_2
X_26359_ _11484_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16112_ _14619_ _14624_ _14525_ VGND VGND VPWR VPWR _14625_ sky130_fd_sc_hd__o21ba_1
XFILLER_196_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29078_ _12952_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__clkbuf_1
X_17092_ _15334_ _15573_ _15576_ _15339_ VGND VGND VPWR VPWR _15577_ sky130_fd_sc_hd__a22o_1
XFILLER_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16043_ _14538_ _14552_ _14554_ _14556_ VGND VGND VPWR VPWR _14557_ sky130_fd_sc_hd__o211a_1
X_28029_ _12395_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31040_ registers\[0\]\[16\] _12968_ _14004_ VGND VGND VPWR VPWR _14011_ sky130_fd_sc_hd__mux2_1
XFILLER_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19802_ _05039_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17994_ _14562_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__buf_6
XFILLER_229_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19733_ registers\[16\]\[38\] registers\[17\]\[38\] registers\[18\]\[38\] registers\[19\]\[38\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16945_ _15434_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32991_ clknet_leaf_42_CLK _01105_ VGND VGND VPWR VPWR registers\[52\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_34730_ clknet_leaf_407_CLK _02844_ VGND VGND VPWR VPWR registers\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_31942_ _09819_ registers\[49\]\[60\] _14418_ VGND VGND VPWR VPWR _14485_ sky130_fd_sc_hd__mux2_1
X_19664_ registers\[20\]\[36\] registers\[21\]\[36\] registers\[22\]\[36\] registers\[23\]\[36\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__mux4_1
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16876_ _15295_ _15366_ _15367_ _15300_ VGND VGND VPWR VPWR _15368_ sky130_fd_sc_hd__a22o_1
XFILLER_226_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18615_ _05122_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__buf_6
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34661_ clknet_leaf_445_CLK _02775_ VGND VGND VPWR VPWR registers\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _06187_ _06322_ _06323_ _06192_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__a22o_1
X_31873_ _09747_ registers\[49\]\[27\] _14441_ VGND VGND VPWR VPWR _14449_ sky130_fd_sc_hd__mux2_1
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33612_ clknet_leaf_171_CLK _01726_ VGND VGND VPWR VPWR registers\[43\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_18546_ _05300_ _05303_ _05074_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__o21ba_1
XFILLER_79_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30824_ _13897_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34592_ clknet_leaf_3_CLK _02706_ VGND VGND VPWR VPWR registers\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33543_ clknet_leaf_255_CLK _01657_ VGND VGND VPWR VPWR registers\[44\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_18477_ registers\[44\]\[3\] registers\[45\]\[3\] registers\[46\]\[3\] registers\[47\]\[3\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__mux4_1
X_30755_ _09676_ registers\[11\]\[9\] _13851_ VGND VGND VPWR VPWR _13861_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_390 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17428_ _14578_ VGND VGND VPWR VPWR _15904_ sky130_fd_sc_hd__buf_4
X_33474_ clknet_leaf_256_CLK _01588_ VGND VGND VPWR VPWR registers\[45\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_30686_ registers\[12\]\[40\] _13018_ _13824_ VGND VGND VPWR VPWR _13825_ sky130_fd_sc_hd__mux2_1
XFILLER_221_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35213_ clknet_leaf_147_CLK _03327_ VGND VGND VPWR VPWR registers\[18\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32425_ clknet_leaf_403_CLK _00539_ VGND VGND VPWR VPWR registers\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36193_ clknet_leaf_29_CLK _00074_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_1
X_17359_ _14592_ VGND VGND VPWR VPWR _15837_ sky130_fd_sc_hd__buf_6
XFILLER_105_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35144_ clknet_leaf_154_CLK _03258_ VGND VGND VPWR VPWR registers\[1\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_20370_ _06919_ _07074_ _07075_ _06922_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__a22o_1
XFILLER_147_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32356_ clknet_leaf_446_CLK _00470_ VGND VGND VPWR VPWR registers\[61\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19029_ registers\[28\]\[18\] registers\[29\]\[18\] registers\[30\]\[18\] registers\[31\]\[18\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__mux4_1
X_31307_ _14151_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__clkbuf_1
X_35075_ clknet_leaf_230_CLK _03189_ VGND VGND VPWR VPWR registers\[20\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32287_ clknet_leaf_2_CLK _00401_ VGND VGND VPWR VPWR registers\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_22040_ _08700_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_8
X_31238_ registers\[8\]\[46\] net41 _14108_ VGND VGND VPWR VPWR _14115_ sky130_fd_sc_hd__mux2_1
XFILLER_115_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34026_ clknet_leaf_426_CLK _02140_ VGND VGND VPWR VPWR registers\[36\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31169_ registers\[8\]\[13\] net5 _14075_ VGND VGND VPWR VPWR _14079_ sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35977_ clknet_leaf_161_CLK _04091_ VGND VGND VPWR VPWR registers\[6\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_23991_ _09531_ registers\[5\]\[8\] _10161_ VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__mux2_1
XFILLER_229_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25730_ _11152_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34928_ clknet_leaf_389_CLK _03042_ VGND VGND VPWR VPWR registers\[22\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_22942_ _09514_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__buf_4
XFILLER_99_1434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25661_ _11116_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22873_ _09487_ _09494_ _09501_ _09508_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__or4_4
X_34859_ clknet_leaf_454_CLK _02973_ VGND VGND VPWR VPWR registers\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_216_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27400_ registers\[36\]\[51\] _10412_ _12062_ VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__mux2_1
XFILLER_227_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24612_ _10529_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28380_ _12580_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__clkbuf_1
X_21824_ _08418_ _08489_ _08490_ _08421_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__a22o_1
X_25592_ _11078_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27331_ _12027_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__clkbuf_1
X_24543_ _10491_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21755_ registers\[28\]\[30\] registers\[29\]\[30\] registers\[30\]\[30\] registers\[31\]\[30\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__mux4_1
XFILLER_51_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20706_ _07276_ _07402_ _07403_ _07286_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__a22o_1
X_27262_ _11935_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__buf_4
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24474_ _10455_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21686_ _08325_ _08340_ _08349_ _08356_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__or4_4
XFILLER_180_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29001_ registers\[24\]\[41\] _10391_ _12905_ VGND VGND VPWR VPWR _12907_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26213_ _10798_ registers\[44\]\[32\] _11405_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__mux2_1
X_23425_ _09654_ _09867_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__nor2_8
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20637_ _07301_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27193_ _11765_ registers\[37\]\[17\] _11947_ VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__mux2_1
XFILLER_137_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26144_ _10729_ _11157_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__nand2_8
XFILLER_137_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23356_ _09831_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
X_20568_ _05107_ _07266_ _07267_ _05117_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__a22o_1
XFILLER_153_915 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22307_ registers\[4\]\[46\] registers\[5\]\[46\] registers\[6\]\[46\] registers\[7\]\[46\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__mux4_1
XFILLER_180_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26075_ _11335_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23287_ registers\[9\]\[45\] _09786_ _09776_ VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__mux2_1
XFILLER_118_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20499_ registers\[8\]\[61\] registers\[9\]\[61\] registers\[10\]\[61\] registers\[11\]\[61\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__mux4_1
XFILLER_124_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29903_ _13412_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__clkbuf_1
X_25026_ net3 VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__buf_2
XFILLER_65_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22238_ registers\[4\]\[44\] registers\[5\]\[44\] registers\[6\]\[44\] registers\[7\]\[44\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__mux4_1
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1706 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1717 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29834_ _13376_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__clkbuf_1
XTAP_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22169_ registers\[0\]\[42\] registers\[1\]\[42\] registers\[2\]\[42\] registers\[3\]\[42\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__mux4_1
XANTENNA_1728 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1739 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29765_ registers\[1\]\[52\] _13044_ _13337_ VGND VGND VPWR VPWR _13340_ sky130_fd_sc_hd__mux2_1
XTAP_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26977_ net46 VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__buf_4
XFILLER_219_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16730_ registers\[20\]\[18\] registers\[21\]\[18\] registers\[22\]\[18\] registers\[23\]\[18\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15226_ sky130_fd_sc_hd__mux4_1
X_28716_ _11801_ registers\[26\]\[34\] _12752_ VGND VGND VPWR VPWR _12757_ sky130_fd_sc_hd__mux2_1
XFILLER_59_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25928_ _10783_ registers\[46\]\[25\] _11252_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__mux2_1
X_29696_ _13303_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16661_ _15129_ _15138_ _15149_ _15158_ VGND VGND VPWR VPWR _15159_ sky130_fd_sc_hd__or4_1
X_25859_ _11221_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
X_28647_ _11732_ registers\[26\]\[1\] _12719_ VGND VGND VPWR VPWR _12721_ sky130_fd_sc_hd__mux2_1
XFILLER_223_919 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18400_ _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16592_ _15091_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
X_19380_ registers\[16\]\[28\] registers\[17\]\[28\] registers\[18\]\[28\] registers\[19\]\[28\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__mux4_1
X_28578_ _12684_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18331_ registers\[60\]\[0\] registers\[61\]\[0\] registers\[62\]\[0\] registers\[63\]\[0\]
+ _05091_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__mux4_1
X_27529_ _12131_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__clkbuf_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18262_ registers\[12\]\[63\] registers\[13\]\[63\] registers\[14\]\[63\] registers\[15\]\[63\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux4_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30540_ _09764_ registers\[13\]\[35\] _13742_ VGND VGND VPWR VPWR _13748_ sky130_fd_sc_hd__mux2_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17213_ _15549_ _15693_ _15694_ _15553_ VGND VGND VPWR VPWR _15695_ sky130_fd_sc_hd__a22o_1
X_30471_ _09662_ registers\[13\]\[2\] _13709_ VGND VGND VPWR VPWR _13712_ sky130_fd_sc_hd__mux2_1
XFILLER_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18193_ registers\[48\]\[61\] registers\[49\]\[61\] registers\[50\]\[61\] registers\[51\]\[61\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__mux4_1
XFILLER_156_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32210_ clknet_leaf_332_CLK _00324_ VGND VGND VPWR VPWR registers\[9\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17144_ registers\[12\]\[30\] registers\[13\]\[30\] registers\[14\]\[30\] registers\[15\]\[30\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15628_ sky130_fd_sc_hd__mux4_1
XFILLER_128_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33190_ clknet_leaf_456_CLK _01304_ VGND VGND VPWR VPWR registers\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32141_ clknet_leaf_460_CLK _00059_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17075_ _14578_ VGND VGND VPWR VPWR _15561_ sky130_fd_sc_hd__buf_4
X_16026_ _14539_ VGND VGND VPWR VPWR _14540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32072_ clknet_leaf_178_CLK _00250_ VGND VGND VPWR VPWR registers\[62\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31023_ registers\[0\]\[8\] _12951_ _13993_ VGND VGND VPWR VPWR _14002_ sky130_fd_sc_hd__mux2_1
X_35900_ clknet_leaf_301_CLK _04014_ VGND VGND VPWR VPWR registers\[7\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35831_ clknet_leaf_318_CLK _03945_ VGND VGND VPWR VPWR registers\[8\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17977_ _04746_ _04749_ _04611_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__o21ba_1
XFILLER_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19716_ _05088_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__clkbuf_4
X_16928_ registers\[8\]\[24\] registers\[9\]\[24\] registers\[10\]\[24\] registers\[11\]\[24\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15418_ sky130_fd_sc_hd__mux4_1
X_35762_ clknet_leaf_382_CLK _03876_ VGND VGND VPWR VPWR registers\[0\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_32974_ clknet_leaf_173_CLK _01088_ VGND VGND VPWR VPWR registers\[52\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34713_ clknet_leaf_20_CLK _02827_ VGND VGND VPWR VPWR registers\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_31925_ _14476_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19647_ _05039_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__buf_4
XFILLER_226_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35693_ clknet_leaf_391_CLK _03807_ VGND VGND VPWR VPWR registers\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16859_ registers\[52\]\[22\] registers\[53\]\[22\] registers\[54\]\[22\] registers\[55\]\[22\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15351_ sky130_fd_sc_hd__mux4_1
XFILLER_93_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34644_ clknet_leaf_93_CLK _02758_ VGND VGND VPWR VPWR registers\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19578_ registers\[52\]\[34\] registers\[53\]\[34\] registers\[54\]\[34\] registers\[55\]\[34\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__mux4_1
X_31856_ _09697_ registers\[49\]\[19\] _14430_ VGND VGND VPWR VPWR _14440_ sky130_fd_sc_hd__mux2_1
XFILLER_240_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18529_ _05111_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__buf_6
X_30807_ _13888_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__clkbuf_1
X_34575_ clknet_leaf_118_CLK _02689_ VGND VGND VPWR VPWR registers\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31787_ registers\[59\]\[50\] net46 _14403_ VGND VGND VPWR VPWR _14404_ sky130_fd_sc_hd__mux2_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33526_ clknet_leaf_340_CLK _01640_ VGND VGND VPWR VPWR registers\[44\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_21540_ registers\[28\]\[24\] registers\[29\]\[24\] registers\[30\]\[24\] registers\[31\]\[24\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__mux4_1
XFILLER_61_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30738_ _13852_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21471_ _08075_ _08146_ _08147_ _08078_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__a22o_1
X_33457_ clknet_leaf_361_CLK _01571_ VGND VGND VPWR VPWR registers\[45\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_30669_ registers\[12\]\[32\] _13002_ _13813_ VGND VGND VPWR VPWR _13816_ sky130_fd_sc_hd__mux2_1
X_23210_ _09736_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_1
X_20422_ _07123_ _07126_ _06880_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__o21ba_1
XFILLER_193_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32408_ clknet_leaf_19_CLK _00522_ VGND VGND VPWR VPWR registers\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_36176_ clknet_leaf_92_CLK _00086_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dfxtp_1
X_24190_ _09594_ registers\[58\]\[38\] _10266_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__mux2_1
XFILLER_162_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33388_ clknet_leaf_345_CLK _01502_ VGND VGND VPWR VPWR registers\[46\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35127_ clknet_leaf_316_CLK _03241_ VGND VGND VPWR VPWR registers\[1\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_23141_ _09694_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
X_20353_ registers\[4\]\[56\] registers\[5\]\[56\] registers\[6\]\[56\] registers\[7\]\[56\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__mux4_1
X_32339_ clknet_leaf_181_CLK _00453_ VGND VGND VPWR VPWR registers\[61\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23072_ _09644_ registers\[62\]\[62\] _09514_ VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__mux2_1
X_20284_ registers\[52\]\[54\] registers\[53\]\[54\] registers\[54\]\[54\] registers\[55\]\[54\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__mux4_1
XFILLER_122_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35058_ clknet_leaf_384_CLK _03172_ VGND VGND VPWR VPWR registers\[20\]\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_11_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_11_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_115_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34009_ clknet_leaf_90_CLK _02123_ VGND VGND VPWR VPWR registers\[36\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_26900_ net18 VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__buf_2
X_22023_ registers\[8\]\[38\] registers\[9\]\[38\] registers\[10\]\[38\] registers\[11\]\[38\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__mux4_1
XTAP_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27880_ _12317_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26831_ _11735_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__clkbuf_1
XTAP_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29550_ registers\[20\]\[14\] _12964_ _13222_ VGND VGND VPWR VPWR _13227_ sky130_fd_sc_hd__mux2_1
XFILLER_57_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26762_ _11697_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_26_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_26_0_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23974_ _10160_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__buf_4
XFILLER_25_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28501_ _12643_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__clkbuf_1
X_25713_ registers\[48\]\[52\] _10414_ _11141_ VGND VGND VPWR VPWR _11144_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22925_ _09545_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
X_26693_ _11661_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_1
X_29481_ _13190_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28432_ _12607_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25644_ _11107_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
X_22856_ registers\[52\]\[63\] registers\[53\]\[63\] registers\[54\]\[63\] registers\[55\]\[63\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__mux4_1
XFILLER_147_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28363_ registers\[2\]\[59\] _10428_ _12561_ VGND VGND VPWR VPWR _12571_ sky130_fd_sc_hd__mux2_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21807_ _08468_ _08473_ _08397_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__o21ba_1
XFILLER_71_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25575_ registers\[4\]\[52\] _10414_ _11067_ VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__mux2_1
XFILLER_169_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22787_ _09148_ _09423_ _09424_ _09153_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__a22o_1
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27314_ registers\[36\]\[10\] _10325_ _12018_ VGND VGND VPWR VPWR _12019_ sky130_fd_sc_hd__mux2_1
XFILLER_80_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24526_ _10482_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28294_ registers\[2\]\[26\] _10359_ _12528_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__mux2_1
X_21738_ _08401_ _08404_ _08405_ _08406_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__o211a_1
XFILLER_160_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27245_ _11982_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_1
X_24457_ _10446_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21669_ _08333_ _08339_ _08062_ _08063_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__o211a_1
XFILLER_184_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23408_ _09858_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27176_ _11748_ registers\[37\]\[9\] _11936_ VGND VGND VPWR VPWR _11946_ sky130_fd_sc_hd__mux2_1
X_24388_ net41 VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26127_ _11362_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
X_23339_ net58 VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__buf_2
X_26058_ _11326_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25009_ _10742_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
X_17900_ _04675_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1503 _07366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18880_ _05350_ _05627_ _05628_ _05353_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__a22o_1
XFILLER_234_1246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1514 _08357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1525 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1536 _09674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17831_ registers\[44\]\[50\] registers\[45\]\[50\] registers\[46\]\[50\] registers\[47\]\[50\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__mux4_1
XANTENNA_1547 _10730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29817_ _13367_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1558 _11585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1569 _12789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17762_ _14531_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__clkbuf_4
X_29748_ registers\[1\]\[44\] _13027_ _13326_ VGND VGND VPWR VPWR _13331_ sky130_fd_sc_hd__mux2_1
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19501_ _06226_ _06229_ _06230_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__a22o_1
XFILLER_169_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16713_ registers\[52\]\[18\] registers\[53\]\[18\] registers\[54\]\[18\] registers\[55\]\[18\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15209_ sky130_fd_sc_hd__mux4_1
XFILLER_208_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17693_ _15884_ _04472_ _04473_ _15890_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__a22o_1
X_29679_ registers\[1\]\[11\] _12958_ _13293_ VGND VGND VPWR VPWR _13295_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_290_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_290_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_169_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31710_ _14363_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__clkbuf_1
X_19432_ _06090_ _06163_ _06164_ _06096_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a22o_1
XFILLER_210_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16644_ _14567_ VGND VGND VPWR VPWR _15142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32690_ clknet_leaf_366_CLK _00804_ VGND VGND VPWR VPWR registers\[57\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31641_ registers\[63\]\[45\] net40 _14321_ VGND VGND VPWR VPWR _14327_ sky130_fd_sc_hd__mux2_1
X_19363_ _05088_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__buf_4
X_16575_ registers\[8\]\[14\] registers\[9\]\[14\] registers\[10\]\[14\] registers\[11\]\[14\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _15075_ sky130_fd_sc_hd__mux4_1
XFILLER_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18314_ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__buf_2
XFILLER_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34360_ clknet_leaf_429_CLK _02474_ VGND VGND VPWR VPWR registers\[31\]\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31572_ registers\[63\]\[12\] net4 _14288_ VGND VGND VPWR VPWR _14291_ sky130_fd_sc_hd__mux2_1
X_19294_ _05039_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__clkbuf_4
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33311_ clknet_leaf_34_CLK _01425_ VGND VGND VPWR VPWR registers\[47\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_18245_ registers\[40\]\[63\] registers\[41\]\[63\] registers\[42\]\[63\] registers\[43\]\[63\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__mux4_1
X_30523_ _09747_ registers\[13\]\[27\] _13731_ VGND VGND VPWR VPWR _13739_ sky130_fd_sc_hd__mux2_1
X_34291_ clknet_leaf_348_CLK _02405_ VGND VGND VPWR VPWR registers\[32\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36030_ clknet_leaf_292_CLK _04144_ VGND VGND VPWR VPWR registers\[63\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_30454_ _13702_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__clkbuf_1
X_33242_ clknet_leaf_35_CLK _01356_ VGND VGND VPWR VPWR registers\[48\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_18176_ registers\[24\]\[60\] registers\[25\]\[60\] registers\[26\]\[60\] registers\[27\]\[60\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__mux4_1
XFILLER_106_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17127_ _15341_ _15609_ _15610_ _15344_ VGND VGND VPWR VPWR _15611_ sky130_fd_sc_hd__a22o_1
XFILLER_89_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33173_ clknet_leaf_78_CLK _01287_ VGND VGND VPWR VPWR registers\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30385_ _13666_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32124_ clknet_leaf_393_CLK _00040_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dfxtp_1
X_17058_ _14541_ VGND VGND VPWR VPWR _15544_ sky130_fd_sc_hd__buf_6
XFILLER_143_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16009_ _14511_ _14514_ _14517_ _14522_ VGND VGND VPWR VPWR _14523_ sky130_fd_sc_hd__a22o_1
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32055_ clknet_leaf_330_CLK _00233_ VGND VGND VPWR VPWR registers\[62\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31006_ _13992_ VGND VGND VPWR VPWR _13993_ sky130_fd_sc_hd__buf_4
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35814_ clknet_leaf_462_CLK _03928_ VGND VGND VPWR VPWR registers\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35745_ clknet_leaf_484_CLK _03859_ VGND VGND VPWR VPWR registers\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_32957_ clknet_leaf_289_CLK _01071_ VGND VGND VPWR VPWR registers\[53\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_20971_ _07586_ _07658_ _07661_ _07589_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_281_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_281_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22710_ registers\[0\]\[58\] registers\[1\]\[58\] registers\[2\]\[58\] registers\[3\]\[58\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__mux4_1
X_31908_ _14467_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__clkbuf_1
X_23690_ registers\[61\]\[60\] _09819_ _09942_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__mux2_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35676_ clknet_leaf_15_CLK _03790_ VGND VGND VPWR VPWR registers\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_32888_ clknet_leaf_331_CLK _01002_ VGND VGND VPWR VPWR registers\[54\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_34627_ clknet_leaf_224_CLK _02741_ VGND VGND VPWR VPWR registers\[27\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_22641_ _09280_ _09283_ _09083_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__o21ba_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31839_ _14431_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25360_ _10764_ registers\[50\]\[16\] _10948_ VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__mux2_1
X_22572_ registers\[32\]\[54\] registers\[33\]\[54\] registers\[34\]\[54\] registers\[35\]\[54\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__mux4_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34558_ clknet_leaf_183_CLK _02672_ VGND VGND VPWR VPWR registers\[28\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24311_ net14 VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__clkbuf_4
XFILLER_221_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33509_ clknet_leaf_59_CLK _01623_ VGND VGND VPWR VPWR registers\[44\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21523_ _07326_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__buf_8
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25291_ _10831_ registers\[51\]\[48\] _10909_ VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__mux2_1
XFILLER_194_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34489_ clknet_leaf_316_CLK _02603_ VGND VGND VPWR VPWR registers\[2\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_27030_ _11869_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36228_ clknet_leaf_121_CLK _00113_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dfxtp_1
X_24242_ _09646_ registers\[58\]\[63\] _10232_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__mux2_1
XFILLER_119_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21454_ _08125_ _08130_ _08054_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__o21ba_1
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20405_ registers\[60\]\[58\] registers\[61\]\[58\] registers\[62\]\[58\] registers\[63\]\[58\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__mux4_1
X_36159_ clknet_leaf_268_CLK _04273_ VGND VGND VPWR VPWR registers\[49\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24173_ _10232_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__clkbuf_8
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21385_ _08058_ _08061_ _08062_ _08063_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__o211a_1
XFILLER_218_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23124_ net4 VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__buf_6
X_20336_ registers\[32\]\[56\] registers\[33\]\[56\] registers\[34\]\[56\] registers\[35\]\[56\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__mux4_1
X_28981_ _12896_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23055_ _09633_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
X_27932_ _12344_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__clkbuf_1
X_20267_ _06873_ _06975_ _06976_ _06878_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__a22o_1
XTAP_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22006_ _08469_ _08665_ _08666_ _08472_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__a22o_1
XTAP_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20198_ _06906_ _06909_ _06880_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__o21ba_1
XTAP_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27863_ _12308_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29602_ registers\[20\]\[39\] _13016_ _13244_ VGND VGND VPWR VPWR _13254_ sky130_fd_sc_hd__mux2_1
XFILLER_236_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26814_ _11724_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__clkbuf_1
XTAP_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27794_ registers\[33\]\[45\] _10399_ _12266_ VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__mux2_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29533_ registers\[20\]\[6\] _12947_ _13211_ VGND VGND VPWR VPWR _13218_ sky130_fd_sc_hd__mux2_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23957_ _10151_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26745_ _11688_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__clkbuf_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_901 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_272_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_272_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22908_ _09533_ registers\[62\]\[9\] _09515_ VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__mux2_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_912 _09708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26676_ _11651_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__clkbuf_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29464_ _13181_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_923 _09802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23888_ _10115_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_934 _10016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_945 _10386_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28415_ _12598_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_956 _10586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22839_ registers\[28\]\[62\] registers\[29\]\[62\] registers\[30\]\[62\] registers\[31\]\[62\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__mux4_1
X_25627_ registers\[48\]\[11\] _10328_ _11097_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__mux2_1
X_29395_ _13145_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_967 _10864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_978 _11229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_989 _11729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16360_ registers\[52\]\[8\] registers\[53\]\[8\] registers\[54\]\[8\] registers\[55\]\[8\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14866_ sky130_fd_sc_hd__mux4_1
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28346_ _12562_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__clkbuf_1
X_25558_ registers\[4\]\[44\] _10397_ _11056_ VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__mux2_1
XFILLER_213_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24509_ _09577_ registers\[56\]\[30\] _10473_ VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__mux2_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16291_ _14567_ VGND VGND VPWR VPWR _14799_ sky130_fd_sc_hd__buf_4
X_28277_ registers\[2\]\[18\] _10342_ _12517_ VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25489_ registers\[4\]\[11\] _10328_ _11023_ VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18030_ registers\[20\]\[55\] registers\[21\]\[55\] registers\[22\]\[55\] registers\[23\]\[55\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__mux4_1
XFILLER_200_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27228_ _11973_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27159_ _11937_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30170_ registers\[16\]\[52\] _13044_ _13550_ VGND VGND VPWR VPWR _13553_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19981_ _06695_ _06698_ _06537_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18932_ registers\[56\]\[16\] registers\[57\]\[16\] registers\[58\]\[16\] registers\[59\]\[16\]
+ _05615_ _05405_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__mux4_1
XANTENNA_1300 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1311 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1322 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1333 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18863_ registers\[36\]\[14\] registers\[37\]\[14\] registers\[38\]\[14\] registers\[39\]\[14\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__mux4_1
XTAP_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1344 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1355 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1366 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17814_ registers\[4\]\[49\] registers\[5\]\[49\] registers\[6\]\[49\] registers\[7\]\[49\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__mux4_1
XANTENNA_1377 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33860_ clknet_leaf_224_CLK _01974_ VGND VGND VPWR VPWR registers\[3\]\[54\] sky130_fd_sc_hd__dfxtp_1
XTAP_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1388 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18794_ _05116_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__clkbuf_4
XTAP_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1399 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32811_ clknet_leaf_422_CLK _00925_ VGND VGND VPWR VPWR registers\[55\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_17745_ registers\[24\]\[47\] registers\[25\]\[47\] registers\[26\]\[47\] registers\[27\]\[47\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__mux4_1
X_33791_ clknet_leaf_273_CLK _01905_ VGND VGND VPWR VPWR registers\[40\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_263_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_263_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35530_ clknet_leaf_151_CLK _03644_ VGND VGND VPWR VPWR registers\[13\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32742_ clknet_leaf_437_CLK _00856_ VGND VGND VPWR VPWR registers\[56\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17676_ registers\[16\]\[45\] registers\[17\]\[45\] registers\[18\]\[45\] registers\[19\]\[45\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__mux4_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19415_ registers\[20\]\[29\] registers\[21\]\[29\] registers\[22\]\[29\] registers\[23\]\[29\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__mux4_1
XFILLER_63_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35461_ clknet_leaf_229_CLK _03575_ VGND VGND VPWR VPWR registers\[14\]\[55\] sky130_fd_sc_hd__dfxtp_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16627_ _14991_ _15123_ _15124_ _14996_ VGND VGND VPWR VPWR _15125_ sky130_fd_sc_hd__a22o_1
XFILLER_223_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32673_ clknet_leaf_43_CLK _00787_ VGND VGND VPWR VPWR registers\[57\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34412_ clknet_leaf_402_CLK _02526_ VGND VGND VPWR VPWR registers\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_31624_ registers\[63\]\[37\] net31 _14310_ VGND VGND VPWR VPWR _14318_ sky130_fd_sc_hd__mux2_1
X_19346_ _06060_ _06067_ _06074_ _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__or4_4
X_35392_ clknet_leaf_238_CLK _03506_ VGND VGND VPWR VPWR registers\[15\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_16558_ _15058_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34343_ clknet_leaf_456_CLK _02457_ VGND VGND VPWR VPWR registers\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31555_ registers\[63\]\[4\] net45 _14277_ VGND VGND VPWR VPWR _14282_ sky130_fd_sc_hd__mux2_1
X_19277_ _06014_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16489_ _14527_ VGND VGND VPWR VPWR _14991_ sky130_fd_sc_hd__clkbuf_4
X_18228_ _04989_ _04992_ _14553_ _14555_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__o211a_1
XFILLER_136_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30506_ _09697_ registers\[13\]\[19\] _13720_ VGND VGND VPWR VPWR _13730_ sky130_fd_sc_hd__mux2_1
XFILLER_248_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34274_ clknet_leaf_48_CLK _02388_ VGND VGND VPWR VPWR registers\[32\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_31486_ _14245_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36013_ clknet_leaf_374_CLK _04127_ VGND VGND VPWR VPWR registers\[63\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_33225_ clknet_leaf_210_CLK _01339_ VGND VGND VPWR VPWR registers\[4\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30437_ _09797_ registers\[14\]\[50\] _13693_ VGND VGND VPWR VPWR _13694_ sky130_fd_sc_hd__mux2_1
X_18159_ registers\[36\]\[60\] registers\[37\]\[60\] registers\[38\]\[60\] registers\[39\]\[60\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux4_1
XFILLER_89_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33156_ clknet_leaf_258_CLK _01270_ VGND VGND VPWR VPWR registers\[50\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21170_ _07326_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__buf_6
XFILLER_137_1206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30368_ _13657_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20121_ registers\[20\]\[49\] registers\[21\]\[49\] registers\[22\]\[49\] registers\[23\]\[49\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux4_1
X_32107_ clknet_leaf_483_CLK _00021_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33087_ clknet_leaf_269_CLK _01201_ VGND VGND VPWR VPWR registers\[51\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_30299_ _13620_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20052_ _06746_ _06753_ _06760_ _06767_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__or4_4
XFILLER_112_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32038_ clknet_leaf_450_CLK _00216_ VGND VGND VPWR VPWR registers\[62\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _09519_ registers\[53\]\[2\] _10658_ VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__mux2_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23811_ _10074_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24791_ _10624_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33989_ clknet_leaf_261_CLK _02103_ VGND VGND VPWR VPWR registers\[37\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_254_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_254_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26530_ _11574_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35728_ clknet_leaf_110_CLK _03842_ VGND VGND VPWR VPWR registers\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_23742_ _09554_ registers\[29\]\[19\] _10028_ VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__mux2_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ registers\[48\]\[8\] registers\[49\]\[8\] registers\[50\]\[8\] registers\[51\]\[8\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__mux4_1
XANTENNA_219 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26461_ _11538_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35659_ clknet_leaf_150_CLK _03773_ VGND VGND VPWR VPWR registers\[11\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_23673_ _10000_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__clkbuf_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ registers\[52\]\[6\] registers\[53\]\[6\] registers\[54\]\[6\] registers\[55\]\[6\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__mux4_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28200_ _12485_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__clkbuf_1
X_25412_ _10982_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
X_22624_ _08958_ _09266_ _09267_ _08961_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__a22o_1
X_29180_ registers\[23\]\[41\] _13021_ _13019_ VGND VGND VPWR VPWR _13022_ sky130_fd_sc_hd__mux2_1
X_26392_ _10842_ registers\[43\]\[53\] _11498_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__mux2_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28131_ _12449_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__clkbuf_1
X_25343_ _10747_ registers\[50\]\[8\] _10937_ VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__mux2_1
XFILLER_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22555_ _08953_ _09199_ _09200_ _08956_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__a22o_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28062_ _11822_ registers\[31\]\[44\] _12408_ VGND VGND VPWR VPWR _12413_ sky130_fd_sc_hd__mux2_1
X_21506_ registers\[28\]\[23\] registers\[29\]\[23\] registers\[30\]\[23\] registers\[31\]\[23\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__mux4_1
XFILLER_195_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25274_ _10864_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__buf_4
X_22486_ registers\[0\]\[51\] registers\[1\]\[51\] registers\[2\]\[51\] registers\[3\]\[51\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__mux4_1
XFILLER_182_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27013_ _11858_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_1
X_24225_ _10293_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
X_21437_ registers\[20\]\[21\] registers\[21\]\[21\] registers\[22\]\[21\] registers\[23\]\[21\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__mux4_1
XFILLER_123_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24156_ _10257_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
X_21368_ registers\[32\]\[20\] registers\[33\]\[20\] registers\[34\]\[20\] registers\[35\]\[20\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__mux4_1
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23107_ _09671_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20319_ registers\[8\]\[55\] registers\[9\]\[55\] registers\[10\]\[55\] registers\[11\]\[55\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__mux4_2
XFILLER_155_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24087_ _10220_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__clkbuf_1
X_28964_ _12887_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__clkbuf_1
X_21299_ registers\[36\]\[18\] registers\[37\]\[18\] registers\[38\]\[18\] registers\[39\]\[18\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__mux4_1
XFILLER_150_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23038_ net47 VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__buf_4
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27915_ _12335_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__clkbuf_1
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28895_ _11845_ registers\[25\]\[55\] _12845_ VGND VGND VPWR VPWR _12851_ sky130_fd_sc_hd__mux2_1
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27846_ _12299_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__clkbuf_1
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27777_ registers\[33\]\[37\] _10382_ _12255_ VGND VGND VPWR VPWR _12263_ sky130_fd_sc_hd__mux2_1
X_24989_ net1 VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__buf_4
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_245_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_245_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29516_ _13208_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__clkbuf_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17530_ _15892_ _04314_ _04315_ _15896_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__a22o_1
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26728_ _11679_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_720 _07340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_731 _07352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_742 _07366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29447_ _13172_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__clkbuf_1
X_17461_ registers\[4\]\[39\] registers\[5\]\[39\] registers\[6\]\[39\] registers\[7\]\[39\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _15936_ sky130_fd_sc_hd__mux4_1
XANTENNA_753 _07385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26659_ _10838_ registers\[41\]\[51\] _11641_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__mux2_1
XFILLER_225_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_764 _07617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_775 _08155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19200_ registers\[4\]\[23\] registers\[5\]\[23\] registers\[6\]\[23\] registers\[7\]\[23\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__mux4_1
XFILLER_220_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16412_ _14895_ _14902_ _14909_ _14916_ VGND VGND VPWR VPWR _14917_ sky130_fd_sc_hd__or4_4
XANTENNA_786 _08804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29378_ _09821_ registers\[22\]\[61\] _13068_ VGND VGND VPWR VPWR _13136_ sky130_fd_sc_hd__mux2_1
XANTENNA_797 _08936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17392_ registers\[24\]\[37\] registers\[25\]\[37\] registers\[26\]\[37\] registers\[27\]\[37\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15869_ sky130_fd_sc_hd__mux4_1
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19131_ _05693_ _05871_ _05872_ _05696_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__a22o_1
X_16343_ registers\[32\]\[8\] registers\[33\]\[8\] registers\[34\]\[8\] registers\[35\]\[8\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14849_ sky130_fd_sc_hd__mux4_1
X_28329_ _12553_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16274_ _14648_ _14780_ _14781_ _14653_ VGND VGND VPWR VPWR _14782_ sky130_fd_sc_hd__a22o_1
XFILLER_200_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19062_ registers\[20\]\[19\] registers\[21\]\[19\] registers\[22\]\[19\] registers\[23\]\[19\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__mux4_1
X_31340_ registers\[7\]\[30\] net24 _14168_ VGND VGND VPWR VPWR _14169_ sky130_fd_sc_hd__mux2_1
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18013_ registers\[48\]\[55\] registers\[49\]\[55\] registers\[50\]\[55\] registers\[51\]\[55\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__mux4_1
XFILLER_172_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31271_ registers\[8\]\[62\] net59 _14063_ VGND VGND VPWR VPWR _14132_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33010_ clknet_leaf_360_CLK _01124_ VGND VGND VPWR VPWR registers\[52\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30222_ _13580_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30153_ registers\[16\]\[44\] _13027_ _13539_ VGND VGND VPWR VPWR _13544_ sky130_fd_sc_hd__mux2_1
X_19964_ _06441_ _06680_ _06681_ _06445_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__a22o_1
XFILLER_214_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18915_ _05659_ _05662_ _05494_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__o21ba_1
XTAP_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34961_ clknet_leaf_114_CLK _03075_ VGND VGND VPWR VPWR registers\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_30084_ registers\[16\]\[11\] _12958_ _13506_ VGND VGND VPWR VPWR _13508_ sky130_fd_sc_hd__mux2_1
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19895_ _06433_ _06613_ _06614_ _06439_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__a22o_1
XANTENNA_1130 _14600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1141 _14667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_484_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_484_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33912_ clknet_leaf_337_CLK _02026_ VGND VGND VPWR VPWR registers\[38\]\[42\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1152 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18846_ registers\[12\]\[13\] registers\[13\]\[13\] registers\[14\]\[13\] registers\[15\]\[13\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__mux4_1
XANTENNA_1163 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34892_ clknet_leaf_144_CLK _03006_ VGND VGND VPWR VPWR registers\[23\]\[62\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1174 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1185 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1196 _15924_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33843_ clknet_leaf_383_CLK _01957_ VGND VGND VPWR VPWR registers\[3\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_18777_ registers\[4\]\[11\] registers\[5\]\[11\] registers\[6\]\[11\] registers\[7\]\[11\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux4_1
X_15989_ _14502_ VGND VGND VPWR VPWR _14503_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_236_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_236_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_208_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17728_ registers\[36\]\[47\] registers\[37\]\[47\] registers\[38\]\[47\] registers\[39\]\[47\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__mux4_1
X_33774_ clknet_leaf_348_CLK _01888_ VGND VGND VPWR VPWR registers\[40\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_30986_ _13982_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35513_ clknet_leaf_303_CLK _03627_ VGND VGND VPWR VPWR registers\[13\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_32725_ clknet_leaf_64_CLK _00839_ VGND VGND VPWR VPWR registers\[56\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17659_ registers\[56\]\[45\] registers\[57\]\[45\] registers\[58\]\[45\] registers\[59\]\[45\]
+ _04408_ _15885_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux4_1
XFILLER_208_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35444_ clknet_leaf_418_CLK _03558_ VGND VGND VPWR VPWR registers\[14\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_20670_ net75 net76 VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__or2_4
X_32656_ clknet_leaf_74_CLK _00770_ VGND VGND VPWR VPWR registers\[57\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19329_ registers\[52\]\[27\] registers\[53\]\[27\] registers\[54\]\[27\] registers\[55\]\[27\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__mux4_1
X_31607_ registers\[63\]\[29\] net22 _14299_ VGND VGND VPWR VPWR _14309_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35375_ clknet_leaf_376_CLK _03489_ VGND VGND VPWR VPWR registers\[15\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32587_ clknet_leaf_150_CLK _00701_ VGND VGND VPWR VPWR registers\[5\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34326_ clknet_leaf_97_CLK _02440_ VGND VGND VPWR VPWR registers\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_22340_ _08953_ _08990_ _08991_ _08956_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__a22o_1
X_31538_ _14272_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34257_ clknet_leaf_132_CLK _02371_ VGND VGND VPWR VPWR registers\[32\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22271_ registers\[12\]\[45\] registers\[13\]\[45\] registers\[14\]\[45\] registers\[15\]\[45\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__mux4_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31469_ _14236_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24010_ _09550_ registers\[5\]\[17\] _10172_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__mux2_1
X_33208_ clknet_leaf_315_CLK _01322_ VGND VGND VPWR VPWR registers\[4\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21222_ _07902_ _07905_ _07744_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__o21ba_1
X_34188_ clknet_leaf_170_CLK _02302_ VGND VGND VPWR VPWR registers\[34\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21153_ registers\[28\]\[13\] registers\[29\]\[13\] registers\[30\]\[13\] registers\[31\]\[13\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__mux4_1
X_33139_ clknet_leaf_364_CLK _01253_ VGND VGND VPWR VPWR registers\[50\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_20104_ registers\[48\]\[49\] registers\[49\]\[49\] registers\[50\]\[49\] registers\[51\]\[49\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__mux4_1
XFILLER_217_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25961_ _11275_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_21084_ registers\[20\]\[11\] registers\[21\]\[11\] registers\[22\]\[11\] registers\[23\]\[11\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__mux4_1
X_27700_ registers\[33\]\[0\] _10303_ _12222_ VGND VGND VPWR VPWR _12223_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_475_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_475_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20035_ registers\[52\]\[47\] registers\[53\]\[47\] registers\[54\]\[47\] registers\[55\]\[47\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__mux4_1
XFILLER_115_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24912_ _09571_ registers\[53\]\[27\] _10680_ VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__mux2_1
X_25892_ _10747_ registers\[46\]\[8\] _11230_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__mux2_1
X_28680_ _11765_ registers\[26\]\[17\] _12730_ VGND VGND VPWR VPWR _12738_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27631_ _12186_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__clkbuf_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24843_ _10651_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_227_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_227_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27562_ _12148_ VGND VGND VPWR VPWR _12149_ sky130_fd_sc_hd__buf_6
X_24774_ _10615_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ registers\[0\]\[37\] registers\[1\]\[37\] registers\[2\]\[37\] registers\[3\]\[37\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__mux4_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_57__f_CLK clknet_5_28_0_CLK VGND VGND VPWR VPWR clknet_6_57__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29301_ _09740_ registers\[22\]\[24\] _13091_ VGND VGND VPWR VPWR _13096_ sky130_fd_sc_hd__mux2_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26513_ _11565_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23725_ _10029_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
X_20937_ registers\[20\]\[7\] registers\[21\]\[7\] registers\[22\]\[7\] registers\[23\]\[7\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__mux4_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27493_ _11795_ registers\[35\]\[31\] _12111_ VGND VGND VPWR VPWR _12113_ sky130_fd_sc_hd__mux2_1
XFILLER_109_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29232_ registers\[23\]\[58\] _13056_ _13040_ VGND VGND VPWR VPWR _13057_ sky130_fd_sc_hd__mux2_1
XFILLER_144_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23656_ _09991_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__clkbuf_1
X_26444_ _11529_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20868_ _07386_ _07560_ _07561_ _07396_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__a22o_1
XFILLER_41_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22607_ _09148_ _09249_ _09250_ _09153_ VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__a22o_1
X_26375_ _10825_ registers\[43\]\[45\] _11487_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__mux2_1
X_29163_ net30 VGND VGND VPWR VPWR _13010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23587_ _09955_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20799_ _07373_ _07493_ _07494_ _07383_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__a22o_1
XFILLER_169_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28114_ _12440_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__clkbuf_1
X_25326_ _10936_ VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22538_ _09184_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29094_ _12963_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25257_ _10900_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__clkbuf_1
X_28045_ _11805_ registers\[31\]\[36\] _12397_ VGND VGND VPWR VPWR _12404_ sky130_fd_sc_hd__mux2_1
X_22469_ _09084_ _09093_ _09103_ _09117_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__or4_4
XFILLER_155_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24208_ _10284_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25188_ _10863_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24139_ _10248_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29996_ _13461_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16961_ _14504_ VGND VGND VPWR VPWR _15450_ sky130_fd_sc_hd__buf_4
X_28947_ _12878_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18700_ _05345_ _05452_ _05453_ _05348_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_466_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_466_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19680_ _06090_ _06404_ _06405_ _06096_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__a22o_1
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28878_ _11828_ registers\[25\]\[47\] _12834_ VGND VGND VPWR VPWR _12842_ sky130_fd_sc_hd__mux2_1
X_16892_ _15206_ _15381_ _15382_ _15210_ VGND VGND VPWR VPWR _15383_ sky130_fd_sc_hd__a22o_1
XFILLER_237_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18631_ _05350_ _05385_ _05386_ _05353_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__a22o_1
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27829_ registers\[33\]\[62\] _10434_ _12221_ VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__mux2_1
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_218_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_218_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18562_ _05316_ _05319_ _05134_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__o21ba_1
X_30840_ _13905_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__clkbuf_1
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17513_ _04294_ _04295_ _04298_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a22o_1
XFILLER_75_1104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ registers\[12\]\[3\] registers\[13\]\[3\] registers\[14\]\[3\] registers\[15\]\[3\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__mux4_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30771_ _13869_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_550 _04539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_561 _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32510_ clknet_leaf_291_CLK _00624_ VGND VGND VPWR VPWR registers\[60\]\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_572 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ registers\[32\]\[39\] registers\[33\]\[39\] registers\[34\]\[39\] registers\[35\]\[39\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _15919_ sky130_fd_sc_hd__mux4_1
X_33490_ clknet_leaf_124_CLK _01604_ VGND VGND VPWR VPWR registers\[44\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_583 _05053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_594 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32441_ clknet_leaf_60_CLK _00555_ VGND VGND VPWR VPWR registers\[29\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17375_ registers\[36\]\[37\] registers\[37\]\[37\] registers\[38\]\[37\] registers\[39\]\[37\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _15852_ sky130_fd_sc_hd__mux4_1
XFILLER_186_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19114_ _05540_ _05854_ _05855_ _05545_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__a22o_1
X_16326_ registers\[8\]\[7\] registers\[9\]\[7\] registers\[10\]\[7\] registers\[11\]\[7\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14833_ sky130_fd_sc_hd__mux4_1
X_35160_ clknet_leaf_8_CLK _03274_ VGND VGND VPWR VPWR registers\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_32372_ clknet_leaf_353_CLK _00486_ VGND VGND VPWR VPWR registers\[61\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34111_ clknet_leaf_269_CLK _02225_ VGND VGND VPWR VPWR registers\[35\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_31323_ registers\[7\]\[22\] net15 _14157_ VGND VGND VPWR VPWR _14160_ sky130_fd_sc_hd__mux2_1
X_19045_ registers\[48\]\[19\] registers\[49\]\[19\] registers\[50\]\[19\] registers\[51\]\[19\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__mux4_1
X_16257_ registers\[0\]\[5\] registers\[1\]\[5\] registers\[2\]\[5\] registers\[3\]\[5\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14766_ sky130_fd_sc_hd__mux4_1
X_35091_ clknet_leaf_105_CLK _03205_ VGND VGND VPWR VPWR registers\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34042_ clknet_leaf_281_CLK _02156_ VGND VGND VPWR VPWR registers\[36\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31254_ _14123_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__clkbuf_1
Xoutput204 net204 VGND VGND VPWR VPWR D2[55] sky130_fd_sc_hd__buf_2
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16188_ registers\[8\]\[3\] registers\[9\]\[3\] registers\[10\]\[3\] registers\[11\]\[3\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _14699_ sky130_fd_sc_hd__mux4_1
Xoutput215 net215 VGND VGND VPWR VPWR D2[7] sky130_fd_sc_hd__buf_2
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput226 net226 VGND VGND VPWR VPWR D3[17] sky130_fd_sc_hd__buf_2
XFILLER_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30205_ _13571_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__clkbuf_1
Xoutput237 net237 VGND VGND VPWR VPWR D3[27] sky130_fd_sc_hd__buf_2
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput248 net248 VGND VGND VPWR VPWR D3[37] sky130_fd_sc_hd__buf_2
XFILLER_86_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput259 net259 VGND VGND VPWR VPWR D3[47] sky130_fd_sc_hd__buf_2
X_31185_ _14087_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19947_ registers\[20\]\[44\] registers\[21\]\[44\] registers\[22\]\[44\] registers\[23\]\[44\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux4_1
X_30136_ registers\[16\]\[36\] _13010_ _13528_ VGND VGND VPWR VPWR _13535_ sky130_fd_sc_hd__mux2_1
XFILLER_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35993_ clknet_leaf_62_CLK _04107_ VGND VGND VPWR VPWR registers\[63\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_457_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_457_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34944_ clknet_leaf_203_CLK _03058_ VGND VGND VPWR VPWR registers\[22\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_30067_ registers\[16\]\[3\] _12941_ _13495_ VGND VGND VPWR VPWR _13499_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19878_ _05125_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__buf_6
XFILLER_114_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ _05540_ _05577_ _05578_ _05545_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a22o_1
X_34875_ clknet_leaf_186_CLK _02989_ VGND VGND VPWR VPWR registers\[23\]\[45\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_209_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_209_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_209_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33826_ clknet_leaf_471_CLK _01940_ VGND VGND VPWR VPWR registers\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_21840_ registers\[56\]\[33\] registers\[57\]\[33\] registers\[58\]\[33\] registers\[59\]\[33\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__mux4_1
XFILLER_243_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21771_ _08435_ _08438_ _08397_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__o21ba_1
X_33757_ clknet_leaf_26_CLK _01871_ VGND VGND VPWR VPWR registers\[40\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_30969_ _13973_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23510_ _09913_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20722_ _07343_ _07418_ _07419_ _07353_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__a22o_1
X_32708_ clknet_leaf_264_CLK _00822_ VGND VGND VPWR VPWR registers\[57\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24490_ _09559_ registers\[56\]\[21\] _10462_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__mux2_1
X_33688_ clknet_leaf_90_CLK _01802_ VGND VGND VPWR VPWR registers\[41\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23441_ _09877_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35427_ clknet_leaf_469_CLK _03541_ VGND VGND VPWR VPWR registers\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_20653_ _07284_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__buf_12
X_32639_ clknet_leaf_268_CLK _00753_ VGND VGND VPWR VPWR registers\[58\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26160_ _10745_ registers\[44\]\[7\] _11372_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__mux2_1
X_35358_ clknet_leaf_484_CLK _03472_ VGND VGND VPWR VPWR registers\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_23372_ _09839_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
X_20584_ registers\[40\]\[0\] registers\[41\]\[0\] registers\[42\]\[0\] registers\[43\]\[0\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__mux4_1
XFILLER_20_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25111_ _10811_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34309_ clknet_leaf_246_CLK _02423_ VGND VGND VPWR VPWR registers\[32\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_22323_ registers\[32\]\[47\] registers\[33\]\[47\] registers\[34\]\[47\] registers\[35\]\[47\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__mux4_1
XFILLER_104_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26091_ _11343_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
X_35289_ clknet_leaf_6_CLK _03403_ VGND VGND VPWR VPWR registers\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25042_ _10764_ registers\[52\]\[16\] _10752_ VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__mux2_1
X_22254_ _08805_ _08906_ _08907_ _08810_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__a22o_1
XFILLER_151_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21205_ _07648_ _07887_ _07888_ _07652_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__a22o_1
X_29850_ _13384_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22185_ _08841_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_2
X_28801_ _11750_ registers\[25\]\[10\] _12801_ VGND VGND VPWR VPWR _12802_ sky130_fd_sc_hd__mux2_1
X_21136_ _07640_ _07820_ _07821_ _07646_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__a22o_1
X_29781_ registers\[1\]\[60\] _13060_ _13281_ VGND VGND VPWR VPWR _13348_ sky130_fd_sc_hd__mux2_1
XFILLER_191_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26993_ net51 VGND VGND VPWR VPWR _11845_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_448_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_448_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_247_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28732_ _12765_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21067_ registers\[48\]\[11\] registers\[49\]\[11\] registers\[50\]\[11\] registers\[51\]\[11\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__mux4_1
X_25944_ _11266_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20018_ _06530_ _06733_ _06734_ _06535_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__a22o_1
X_28663_ _11748_ registers\[26\]\[9\] _12719_ VGND VGND VPWR VPWR _12729_ sky130_fd_sc_hd__mux2_1
X_25875_ _11229_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__buf_4
XFILLER_150_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27614_ _12177_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__clkbuf_1
X_24826_ _09619_ registers\[54\]\[50\] _10642_ VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__mux2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28594_ _11813_ registers\[27\]\[40\] _12692_ VGND VGND VPWR VPWR _12693_ sky130_fd_sc_hd__mux2_1
XFILLER_64_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27545_ _11847_ registers\[35\]\[56\] _12133_ VGND VGND VPWR VPWR _12140_ sky130_fd_sc_hd__mux2_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ registers\[40\]\[37\] registers\[41\]\[37\] registers\[42\]\[37\] registers\[43\]\[37\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__mux4_1
XFILLER_76_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24757_ _10606_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23708_ _10020_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkbuf_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24688_ _10513_ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__clkbuf_8
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27476_ _11778_ registers\[35\]\[23\] _12100_ VGND VGND VPWR VPWR _12104_ sky130_fd_sc_hd__mux2_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29215_ _13045_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26427_ _11520_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__clkbuf_1
X_23639_ _09982_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__clkbuf_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_773 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29146_ registers\[23\]\[30\] _12997_ _12998_ VGND VGND VPWR VPWR _12999_ sky130_fd_sc_hd__mux2_1
X_17160_ _15638_ _15639_ _15642_ _15643_ VGND VGND VPWR VPWR _15644_ sky130_fd_sc_hd__a22o_1
XFILLER_211_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26358_ _10808_ registers\[43\]\[37\] _11476_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__mux2_1
XFILLER_156_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16111_ _14511_ _14620_ _14623_ _14517_ VGND VGND VPWR VPWR _14624_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25309_ _10927_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_1
X_26289_ _10739_ registers\[43\]\[4\] _11443_ VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__mux2_1
X_29077_ registers\[23\]\[8\] _12951_ _12935_ VGND VGND VPWR VPWR _12952_ sky130_fd_sc_hd__mux2_1
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17091_ registers\[32\]\[29\] registers\[33\]\[29\] registers\[34\]\[29\] registers\[35\]\[29\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15576_ sky130_fd_sc_hd__mux4_1
XFILLER_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16042_ _14555_ VGND VGND VPWR VPWR _14556_ sky130_fd_sc_hd__buf_2
X_28028_ _11788_ registers\[31\]\[28\] _12386_ VGND VGND VPWR VPWR _12395_ sky130_fd_sc_hd__mux2_1
XFILLER_124_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19801_ _06519_ _06522_ _06523_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__o21ba_1
XFILLER_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17993_ _04762_ _04765_ _04630_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__o21ba_1
X_29979_ _13452_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_439_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_439_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19732_ registers\[24\]\[38\] registers\[25\]\[38\] registers\[26\]\[38\] registers\[27\]\[38\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__mux4_1
XFILLER_42_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16944_ _15408_ _15417_ _15424_ _15433_ VGND VGND VPWR VPWR _15434_ sky130_fd_sc_hd__or4_4
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32990_ clknet_leaf_42_CLK _01104_ VGND VGND VPWR VPWR registers\[52\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31941_ _14484_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19663_ registers\[28\]\[36\] registers\[29\]\[36\] registers\[30\]\[36\] registers\[31\]\[36\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__mux4_1
X_16875_ registers\[20\]\[22\] registers\[21\]\[22\] registers\[22\]\[22\] registers\[23\]\[22\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15367_ sky130_fd_sc_hd__mux4_1
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18614_ _05120_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__buf_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34660_ clknet_leaf_474_CLK _02774_ VGND VGND VPWR VPWR registers\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ registers\[20\]\[34\] registers\[21\]\[34\] registers\[22\]\[34\] registers\[23\]\[34\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__mux4_1
X_31872_ _14448_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33611_ clknet_leaf_159_CLK _01725_ VGND VGND VPWR VPWR registers\[43\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_18545_ _05204_ _05301_ _05302_ _05207_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__a22o_1
XFILLER_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30823_ _09778_ registers\[11\]\[41\] _13895_ VGND VGND VPWR VPWR _13897_ sky130_fd_sc_hd__mux2_1
X_34591_ clknet_leaf_9_CLK _02705_ VGND VGND VPWR VPWR registers\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_40__f_CLK clknet_5_20_0_CLK VGND VGND VPWR VPWR clknet_6_40__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_234_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33542_ clknet_leaf_254_CLK _01656_ VGND VGND VPWR VPWR registers\[44\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_18476_ _05197_ _05234_ _05235_ _05202_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__a22o_1
X_30754_ _13860_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_863 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_380 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_391 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ _14576_ VGND VGND VPWR VPWR _15903_ sky130_fd_sc_hd__buf_6
X_33473_ clknet_leaf_257_CLK _01587_ VGND VGND VPWR VPWR registers\[45\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30685_ _13779_ VGND VGND VPWR VPWR _13824_ sky130_fd_sc_hd__buf_4
XFILLER_92_1292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35212_ clknet_leaf_147_CLK _03326_ VGND VGND VPWR VPWR registers\[18\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32424_ clknet_leaf_454_CLK _00538_ VGND VGND VPWR VPWR registers\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_36192_ clknet_leaf_29_CLK _00073_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_1
X_17358_ registers\[24\]\[36\] registers\[25\]\[36\] registers\[26\]\[36\] registers\[27\]\[36\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15836_ sky130_fd_sc_hd__mux4_1
XFILLER_118_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35143_ clknet_leaf_154_CLK _03257_ VGND VGND VPWR VPWR registers\[1\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_16309_ _14816_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
X_32355_ clknet_leaf_445_CLK _00469_ VGND VGND VPWR VPWR registers\[61\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17289_ _14564_ VGND VGND VPWR VPWR _15769_ sky130_fd_sc_hd__buf_4
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19028_ _05496_ _05771_ _05772_ _05499_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a22o_1
X_31306_ registers\[7\]\[14\] net6 _14146_ VGND VGND VPWR VPWR _14151_ sky130_fd_sc_hd__mux2_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35074_ clknet_leaf_230_CLK _03188_ VGND VGND VPWR VPWR registers\[20\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_32286_ clknet_leaf_3_CLK _00400_ VGND VGND VPWR VPWR registers\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_34025_ clknet_leaf_425_CLK _02139_ VGND VGND VPWR VPWR registers\[36\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31237_ _14114_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31168_ _14078_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30119_ registers\[16\]\[28\] _12993_ _13517_ VGND VGND VPWR VPWR _13526_ sky130_fd_sc_hd__mux2_1
X_23990_ _10169_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35976_ clknet_leaf_160_CLK _04090_ VGND VGND VPWR VPWR registers\[6\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31099_ registers\[0\]\[44\] _13027_ _14037_ VGND VGND VPWR VPWR _14042_ sky130_fd_sc_hd__mux2_1
XFILLER_229_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22941_ net13 VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__buf_2
XFILLER_214_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34927_ clknet_leaf_387_CLK _03041_ VGND VGND VPWR VPWR registers\[22\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22872_ _09504_ _09507_ _07398_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__o21ba_1
XFILLER_216_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25660_ registers\[48\]\[27\] _10361_ _11108_ VGND VGND VPWR VPWR _11116_ sky130_fd_sc_hd__mux2_1
XFILLER_228_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34858_ clknet_leaf_453_CLK _02972_ VGND VGND VPWR VPWR registers\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24611_ _09542_ registers\[55\]\[13\] _10525_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__mux2_1
X_21823_ registers\[16\]\[32\] registers\[17\]\[32\] registers\[18\]\[32\] registers\[19\]\[32\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__mux4_1
X_25591_ registers\[4\]\[60\] _10430_ _11011_ VGND VGND VPWR VPWR _11078_ sky130_fd_sc_hd__mux2_1
X_33809_ clknet_leaf_109_CLK _01923_ VGND VGND VPWR VPWR registers\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34789_ clknet_leaf_446_CLK _02903_ VGND VGND VPWR VPWR registers\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24542_ _09611_ registers\[56\]\[46\] _10484_ VGND VGND VPWR VPWR _10491_ sky130_fd_sc_hd__mux2_1
X_27330_ registers\[36\]\[18\] _10342_ _12018_ VGND VGND VPWR VPWR _12027_ sky130_fd_sc_hd__mux2_1
X_21754_ _07385_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20705_ registers\[32\]\[1\] registers\[33\]\[1\] registers\[34\]\[1\] registers\[35\]\[1\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__mux4_1
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27261_ _11990_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24473_ _09542_ registers\[56\]\[13\] _10451_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__mux2_1
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21685_ _08352_ _08355_ _08087_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__o21ba_1
XFILLER_225_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29000_ _12906_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23424_ net85 net84 VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__nand2b_4
X_26212_ _11407_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
X_20636_ registers\[52\]\[0\] registers\[53\]\[0\] registers\[54\]\[0\] registers\[55\]\[0\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__mux4_1
X_27192_ _11954_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26143_ _11370_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23355_ registers\[39\]\[31\] _09756_ _09829_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__mux2_1
X_20567_ registers\[16\]\[63\] registers\[17\]\[63\] registers\[18\]\[63\] registers\[19\]\[63\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__mux4_1
XFILLER_50_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22306_ registers\[12\]\[46\] registers\[13\]\[46\] registers\[14\]\[46\] registers\[15\]\[46\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__mux4_1
X_26074_ _10793_ registers\[45\]\[30\] _11334_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23286_ net40 VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__clkbuf_4
X_20498_ _07196_ _07199_ _05102_ _05104_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__o211a_1
XFILLER_180_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29902_ registers\[18\]\[53\] _13046_ _13408_ VGND VGND VPWR VPWR _13412_ sky130_fd_sc_hd__mux2_1
X_25025_ _10753_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22237_ registers\[12\]\[44\] registers\[13\]\[44\] registers\[14\]\[44\] registers\[15\]\[44\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__mux4_1
XFILLER_65_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29833_ registers\[18\]\[20\] _12976_ _13375_ VGND VGND VPWR VPWR _13376_ sky130_fd_sc_hd__mux2_1
XANTENNA_1707 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22168_ registers\[8\]\[42\] registers\[9\]\[42\] registers\[10\]\[42\] registers\[11\]\[42\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__mux4_1
XTAP_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1718 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1729 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21119_ _07377_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__buf_6
XTAP_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29764_ _13339_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26976_ _11833_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22099_ _08615_ _08756_ _08757_ _08618_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__a22o_1
XTAP_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28715_ _12756_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25927_ _11257_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
X_29695_ registers\[1\]\[19\] _12974_ _13293_ VGND VGND VPWR VPWR _13303_ sky130_fd_sc_hd__mux2_1
XFILLER_75_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28646_ _12720_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16660_ _15154_ _15157_ _14959_ VGND VGND VPWR VPWR _15158_ sky130_fd_sc_hd__o21ba_1
X_25858_ _10848_ registers\[47\]\[56\] _11214_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24809_ _09603_ registers\[54\]\[42\] _10631_ VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__mux2_1
X_28577_ _11797_ registers\[27\]\[32\] _12681_ VGND VGND VPWR VPWR _12684_ sky130_fd_sc_hd__mux2_1
X_16591_ _15065_ _15074_ _15081_ _15090_ VGND VGND VPWR VPWR _15091_ sky130_fd_sc_hd__or4_1
XFILLER_222_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25789_ _10779_ registers\[47\]\[23\] _11181_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__mux2_1
XFILLER_243_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18330_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__buf_4
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27528_ _11830_ registers\[35\]\[48\] _12122_ VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__mux2_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _14491_ _05023_ _05024_ _14501_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__a22o_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27459_ _11761_ registers\[35\]\[15\] _12089_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__mux2_1
XFILLER_230_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17212_ registers\[52\]\[32\] registers\[53\]\[32\] registers\[54\]\[32\] registers\[55\]\[32\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15694_ sky130_fd_sc_hd__mux4_1
XFILLER_243_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30470_ _13711_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__clkbuf_1
X_18192_ registers\[56\]\[61\] registers\[57\]\[61\] registers\[58\]\[61\] registers\[59\]\[61\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__mux4_1
XFILLER_168_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17143_ _15482_ _15623_ _15626_ _15485_ VGND VGND VPWR VPWR _15627_ sky130_fd_sc_hd__a22o_1
X_29129_ net18 VGND VGND VPWR VPWR _12987_ sky130_fd_sc_hd__buf_2
XFILLER_11_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32140_ clknet_leaf_462_CLK _00058_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17074_ _14576_ VGND VGND VPWR VPWR _15560_ sky130_fd_sc_hd__buf_6
XFILLER_155_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16025_ _14509_ VGND VGND VPWR VPWR _14539_ sky130_fd_sc_hd__buf_12
X_32071_ clknet_leaf_195_CLK _00249_ VGND VGND VPWR VPWR registers\[62\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31022_ _14001_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35830_ clknet_leaf_330_CLK _03944_ VGND VGND VPWR VPWR registers\[8\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_17976_ _04683_ _04747_ _04748_ _04686_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__a22o_1
XFILLER_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19715_ _06433_ _06435_ _06438_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__a22o_1
XFILLER_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16927_ _15412_ _15416_ _15277_ _15278_ VGND VGND VPWR VPWR _15417_ sky130_fd_sc_hd__o211a_1
XFILLER_66_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32973_ clknet_leaf_142_CLK _01087_ VGND VGND VPWR VPWR registers\[53\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_35761_ clknet_leaf_381_CLK _03875_ VGND VGND VPWR VPWR registers\[0\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31924_ _09800_ registers\[49\]\[51\] _14474_ VGND VGND VPWR VPWR _14476_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19646_ _06367_ _06372_ _06169_ _06170_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__o211a_1
X_34712_ clknet_leaf_18_CLK _02826_ VGND VGND VPWR VPWR registers\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35692_ clknet_leaf_392_CLK _03806_ VGND VGND VPWR VPWR registers\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_16858_ registers\[60\]\[22\] registers\[61\]\[22\] registers\[62\]\[22\] registers\[63\]\[22\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15350_ sky130_fd_sc_hd__mux4_1
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34643_ clknet_leaf_104_CLK _02757_ VGND VGND VPWR VPWR registers\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19577_ registers\[60\]\[34\] registers\[61\]\[34\] registers\[62\]\[34\] registers\[63\]\[34\]
+ _06305_ _06099_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__mux4_1
XFILLER_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31855_ _14439_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16789_ registers\[0\]\[20\] registers\[1\]\[20\] registers\[2\]\[20\] registers\[3\]\[20\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15283_ sky130_fd_sc_hd__mux4_1
XFILLER_225_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18528_ _05283_ _05286_ _05134_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__o21ba_1
X_30806_ _09760_ registers\[11\]\[33\] _13884_ VGND VGND VPWR VPWR _13888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34574_ clknet_leaf_119_CLK _02688_ VGND VGND VPWR VPWR registers\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_31786_ _14347_ VGND VGND VPWR VPWR _14403_ sky130_fd_sc_hd__buf_6
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33525_ clknet_leaf_345_CLK _01639_ VGND VGND VPWR VPWR registers\[44\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_18459_ registers\[12\]\[2\] registers\[13\]\[2\] registers\[14\]\[2\] registers\[15\]\[2\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__mux4_1
X_30737_ _09648_ registers\[11\]\[0\] _13851_ VGND VGND VPWR VPWR _13852_ sky130_fd_sc_hd__mux2_1
XFILLER_194_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33456_ clknet_leaf_362_CLK _01570_ VGND VGND VPWR VPWR registers\[45\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_21470_ registers\[16\]\[22\] registers\[17\]\[22\] registers\[18\]\[22\] registers\[19\]\[22\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__mux4_1
X_30668_ _13815_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20421_ _06873_ _07124_ _07125_ _06878_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__a22o_1
X_32407_ clknet_leaf_93_CLK _00521_ VGND VGND VPWR VPWR registers\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_36175_ clknet_leaf_92_CLK _00075_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33387_ clknet_leaf_429_CLK _01501_ VGND VGND VPWR VPWR registers\[46\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_30599_ _13778_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35126_ clknet_leaf_317_CLK _03240_ VGND VGND VPWR VPWR registers\[1\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_23140_ registers\[39\]\[17\] _09693_ _09679_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__mux2_1
X_20352_ registers\[12\]\[56\] registers\[13\]\[56\] registers\[14\]\[56\] registers\[15\]\[56\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__mux4_1
X_32338_ clknet_leaf_72_CLK _00452_ VGND VGND VPWR VPWR registers\[61\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23071_ net59 VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__buf_2
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35057_ clknet_leaf_385_CLK _03171_ VGND VGND VPWR VPWR registers\[20\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_32269_ clknet_leaf_168_CLK _00383_ VGND VGND VPWR VPWR registers\[39\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20283_ registers\[60\]\[54\] registers\[61\]\[54\] registers\[62\]\[54\] registers\[63\]\[54\]
+ _06991_ _06785_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__mux4_1
XFILLER_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34008_ clknet_leaf_90_CLK _02122_ VGND VGND VPWR VPWR registers\[36\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_22022_ _08676_ _08682_ _08405_ _08406_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__o211a_1
XTAP_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26830_ _11734_ registers\[3\]\[2\] _11730_ VGND VGND VPWR VPWR _11735_ sky130_fd_sc_hd__mux2_1
XTAP_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26761_ registers\[40\]\[35\] _10378_ _11691_ VGND VGND VPWR VPWR _11697_ sky130_fd_sc_hd__mux2_1
X_23973_ _10015_ _10159_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__nand2_8
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35959_ clknet_leaf_313_CLK _04073_ VGND VGND VPWR VPWR registers\[6\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28500_ _11855_ registers\[28\]\[60\] _12576_ VGND VGND VPWR VPWR _12643_ sky130_fd_sc_hd__mux2_1
X_25712_ _11143_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29480_ _09786_ registers\[21\]\[45\] _13184_ VGND VGND VPWR VPWR _13190_ sky130_fd_sc_hd__mux2_1
X_22924_ _09544_ registers\[62\]\[14\] _09536_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__mux2_1
XFILLER_244_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26692_ registers\[40\]\[2\] _10309_ _11658_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28431_ _11786_ registers\[28\]\[27\] _12599_ VGND VGND VPWR VPWR _12607_ sky130_fd_sc_hd__mux2_1
XFILLER_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25643_ registers\[48\]\[19\] _10344_ _11097_ VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__mux2_1
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22855_ registers\[60\]\[63\] registers\[61\]\[63\] registers\[62\]\[63\] registers\[63\]\[63\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__mux4_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28362_ _12570_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_1
X_21806_ _08469_ _08470_ _08471_ _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__a22o_1
XFILLER_73_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22786_ registers\[32\]\[61\] registers\[33\]\[61\] registers\[34\]\[61\] registers\[35\]\[61\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__mux4_1
XFILLER_213_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25574_ _11069_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27313_ _12006_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__buf_4
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21737_ _07340_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__clkbuf_4
X_24525_ _09594_ registers\[56\]\[38\] _10473_ VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__mux2_1
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28293_ _12534_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27244_ _11816_ registers\[37\]\[41\] _11980_ VGND VGND VPWR VPWR _11982_ sky130_fd_sc_hd__mux2_1
X_24456_ _09525_ registers\[56\]\[5\] _10440_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__mux2_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21668_ _08334_ _08336_ _08337_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__a22o_1
XFILLER_123_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23407_ registers\[39\]\[56\] _09810_ _09851_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__mux2_1
X_20619_ registers\[56\]\[0\] registers\[57\]\[0\] registers\[58\]\[0\] registers\[59\]\[0\]
+ _07315_ _07317_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__mux4_1
X_27175_ _11945_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__clkbuf_1
X_24387_ _10400_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21599_ _07295_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__clkbuf_4
X_23338_ _09820_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
X_26126_ _10846_ registers\[45\]\[55\] _11356_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__mux2_1
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26057_ _10777_ registers\[45\]\[22\] _11323_ VGND VGND VPWR VPWR _11326_ sky130_fd_sc_hd__mux2_1
X_23269_ _09774_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_4__f_CLK clknet_5_2_0_CLK VGND VGND VPWR VPWR clknet_6_4__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25008_ _10741_ registers\[52\]\[5\] _10731_ VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__mux2_1
XFILLER_152_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1504 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1515 _08357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1526 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ _14548_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__clkbuf_4
X_29816_ registers\[18\]\[12\] _12960_ _13364_ VGND VGND VPWR VPWR _13367_ sky130_fd_sc_hd__mux2_1
XTAP_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1537 _09780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1548 _10730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1559 _11585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _14489_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29747_ _13330_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__clkbuf_1
X_26959_ net39 VGND VGND VPWR VPWR _11822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19500_ _05049_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__buf_2
X_16712_ registers\[60\]\[18\] registers\[61\]\[18\] registers\[62\]\[18\] registers\[63\]\[18\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15208_ sky130_fd_sc_hd__mux4_1
XFILLER_43_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17692_ registers\[48\]\[46\] registers\[49\]\[46\] registers\[50\]\[46\] registers\[51\]\[46\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__mux4_1
X_29678_ _13294_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19431_ registers\[48\]\[30\] registers\[49\]\[30\] registers\[50\]\[30\] registers\[51\]\[30\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__mux4_1
X_28629_ _11849_ registers\[27\]\[57\] _12703_ VGND VGND VPWR VPWR _12711_ sky130_fd_sc_hd__mux2_1
X_16643_ registers\[0\]\[16\] registers\[1\]\[16\] registers\[2\]\[16\] registers\[3\]\[16\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15141_ sky130_fd_sc_hd__mux4_1
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31640_ _14326_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__clkbuf_1
X_19362_ _06090_ _06092_ _06095_ _06096_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__a22o_1
X_16574_ _15069_ _15073_ _14934_ _14935_ VGND VGND VPWR VPWR _15074_ sky130_fd_sc_hd__o211a_2
XFILLER_231_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18313_ _05038_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__buf_12
XFILLER_163_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31571_ _14290_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__clkbuf_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19293_ _06024_ _06029_ _05826_ _05827_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__o211a_1
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33310_ clknet_leaf_28_CLK _01424_ VGND VGND VPWR VPWR registers\[47\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_18244_ _05008_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
X_30522_ _13738_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__clkbuf_1
X_34290_ clknet_leaf_360_CLK _02404_ VGND VGND VPWR VPWR registers\[32\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33241_ clknet_leaf_35_CLK _01355_ VGND VGND VPWR VPWR registers\[48\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18175_ _04938_ _04941_ _14584_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__o21ba_1
X_30453_ _09815_ registers\[14\]\[58\] _13693_ VGND VGND VPWR VPWR _13702_ sky130_fd_sc_hd__mux2_1
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17126_ registers\[36\]\[30\] registers\[37\]\[30\] registers\[38\]\[30\] registers\[39\]\[30\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15610_ sky130_fd_sc_hd__mux4_1
X_33172_ clknet_leaf_70_CLK _01286_ VGND VGND VPWR VPWR registers\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_30384_ _09742_ registers\[14\]\[25\] _13660_ VGND VGND VPWR VPWR _13666_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32123_ clknet_leaf_397_CLK _00039_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dfxtp_1
X_17057_ registers\[56\]\[28\] registers\[57\]\[28\] registers\[58\]\[28\] registers\[59\]\[28\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15543_ sky130_fd_sc_hd__mux4_1
XFILLER_83_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16008_ registers\[36\]\[0\] registers\[37\]\[0\] registers\[38\]\[0\] registers\[39\]\[0\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14522_ sky130_fd_sc_hd__mux4_1
XFILLER_143_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32054_ clknet_leaf_330_CLK _00232_ VGND VGND VPWR VPWR registers\[62\]\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31005_ _11008_ _11084_ VGND VGND VPWR VPWR _13992_ sky130_fd_sc_hd__nor2_8
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35813_ clknet_leaf_462_CLK _03927_ VGND VGND VPWR VPWR registers\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17959_ registers\[4\]\[53\] registers\[5\]\[53\] registers\[6\]\[53\] registers\[7\]\[53\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux4_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32956_ clknet_leaf_290_CLK _01070_ VGND VGND VPWR VPWR registers\[53\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_20970_ registers\[4\]\[8\] registers\[5\]\[8\] registers\[6\]\[8\] registers\[7\]\[8\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__mux4_1
X_35744_ clknet_leaf_486_CLK _03858_ VGND VGND VPWR VPWR registers\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31907_ _09782_ registers\[49\]\[43\] _14463_ VGND VGND VPWR VPWR _14467_ sky130_fd_sc_hd__mux2_1
X_19629_ _06333_ _06340_ _06349_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__or4_1
X_35675_ clknet_leaf_14_CLK _03789_ VGND VGND VPWR VPWR registers\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_32887_ clknet_leaf_330_CLK _01001_ VGND VGND VPWR VPWR registers\[54\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_22640_ _09155_ _09281_ _09282_ _09158_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__a22o_1
XFILLER_81_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34626_ clknet_leaf_224_CLK _02740_ VGND VGND VPWR VPWR registers\[27\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_31838_ _09678_ registers\[49\]\[10\] _14430_ VGND VGND VPWR VPWR _14431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22571_ registers\[40\]\[54\] registers\[41\]\[54\] registers\[42\]\[54\] registers\[43\]\[54\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__mux4_1
X_34557_ clknet_leaf_183_CLK _02671_ VGND VGND VPWR VPWR registers\[28\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31769_ _14394_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24310_ _10348_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
X_21522_ _07983_ _08195_ _08196_ _07989_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__a22o_1
X_25290_ _10917_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__clkbuf_1
X_33508_ clknet_leaf_61_CLK _01622_ VGND VGND VPWR VPWR registers\[44\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34488_ clknet_leaf_316_CLK _02602_ VGND VGND VPWR VPWR registers\[2\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24241_ _10301_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36227_ clknet_leaf_121_CLK _00112_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dfxtp_1
X_21453_ _08126_ _08127_ _08128_ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__a22o_1
X_33439_ clknet_leaf_33_CLK _01553_ VGND VGND VPWR VPWR registers\[45\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20404_ _05136_ _07107_ _07108_ _05146_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__a22o_1
XFILLER_193_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36158_ clknet_leaf_268_CLK _04272_ VGND VGND VPWR VPWR registers\[49\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24172_ _10265_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21384_ _07340_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__clkbuf_4
X_23123_ _09682_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
X_20335_ registers\[40\]\[56\] registers\[41\]\[56\] registers\[42\]\[56\] registers\[43\]\[56\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__mux4_1
X_35109_ clknet_leaf_465_CLK _03223_ VGND VGND VPWR VPWR registers\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36089_ clknet_leaf_333_CLK _04203_ VGND VGND VPWR VPWR registers\[59\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_28980_ registers\[24\]\[31\] _10370_ _12894_ VGND VGND VPWR VPWR _12896_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23054_ _09632_ registers\[62\]\[56\] _09620_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__mux2_1
X_27931_ registers\[32\]\[46\] _10401_ _12337_ VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__mux2_1
X_20266_ registers\[20\]\[53\] registers\[21\]\[53\] registers\[22\]\[53\] registers\[23\]\[53\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__mux4_1
XTAP_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22005_ registers\[36\]\[38\] registers\[37\]\[38\] registers\[38\]\[38\] registers\[39\]\[38\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__mux4_1
XTAP_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27862_ registers\[32\]\[13\] _10332_ _12304_ VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__mux2_1
X_20197_ _06873_ _06907_ _06908_ _06878_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__a22o_1
XTAP_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29601_ _13253_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26813_ registers\[40\]\[60\] _10430_ _11657_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__mux2_1
XTAP_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27793_ _12271_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__clkbuf_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29532_ _13217_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__clkbuf_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26744_ registers\[40\]\[27\] _10361_ _11680_ VGND VGND VPWR VPWR _11688_ sky130_fd_sc_hd__mux2_1
X_23956_ _09632_ registers\[60\]\[56\] _10144_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__mux2_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1010 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_902 _09660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22907_ net64 VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__clkbuf_4
X_29463_ _09769_ registers\[21\]\[37\] _13173_ VGND VGND VPWR VPWR _13181_ sky130_fd_sc_hd__mux2_1
X_26675_ _10854_ registers\[41\]\[59\] _11641_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_913 _09708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_924 _09810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _09563_ registers\[60\]\[23\] _10111_ VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_935 _10160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28414_ _11769_ registers\[28\]\[19\] _12588_ VGND VGND VPWR VPWR _12598_ sky130_fd_sc_hd__mux2_1
X_25626_ _11098_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_946 _10391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22838_ _07343_ _09473_ _09474_ _07353_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__a22o_1
X_29394_ _09666_ registers\[21\]\[4\] _13140_ VGND VGND VPWR VPWR _13145_ sky130_fd_sc_hd__mux2_1
XANTENNA_957 _10586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_968 _10936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_979 _11229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28345_ registers\[2\]\[50\] _10409_ _12561_ VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__mux2_1
XFILLER_227_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25557_ _11060_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__clkbuf_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22769_ registers\[8\]\[60\] registers\[9\]\[60\] registers\[10\]\[60\] registers\[11\]\[60\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__mux4_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24508_ _10439_ VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__clkbuf_8
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ registers\[0\]\[6\] registers\[1\]\[6\] registers\[2\]\[6\] registers\[3\]\[6\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14798_ sky130_fd_sc_hd__mux4_1
X_28276_ _12525_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__clkbuf_1
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25488_ _11024_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27227_ _11799_ registers\[37\]\[33\] _11969_ VGND VGND VPWR VPWR _11973_ sky130_fd_sc_hd__mux2_1
X_24439_ _10435_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
X_27158_ _11728_ registers\[37\]\[0\] _11936_ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__mux2_1
X_26109_ _10829_ registers\[45\]\[47\] _11345_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__mux2_1
X_19980_ _06530_ _06696_ _06697_ _06535_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__a22o_1
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27089_ _11900_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18931_ _05674_ _05677_ _05475_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__o21ba_1
XFILLER_234_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1301 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1312 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1323 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18862_ registers\[44\]\[14\] registers\[45\]\[14\] registers\[46\]\[14\] registers\[47\]\[14\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__mux4_1
XTAP_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1334 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1345 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17813_ registers\[12\]\[49\] registers\[13\]\[49\] registers\[14\]\[49\] registers\[15\]\[49\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__mux4_1
XFILLER_67_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1356 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1367 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1378 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18793_ registers\[32\]\[12\] registers\[33\]\[12\] registers\[34\]\[12\] registers\[35\]\[12\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__mux4_1
XTAP_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1389 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_212_1342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32810_ clknet_leaf_422_CLK _00924_ VGND VGND VPWR VPWR registers\[55\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ _04520_ _04523_ _15974_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__o21ba_1
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33790_ clknet_leaf_273_CLK _01904_ VGND VGND VPWR VPWR registers\[40\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32741_ clknet_leaf_438_CLK _00855_ VGND VGND VPWR VPWR registers\[56\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_17675_ registers\[24\]\[45\] registers\[25\]\[45\] registers\[26\]\[45\] registers\[27\]\[45\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19414_ registers\[28\]\[29\] registers\[29\]\[29\] registers\[30\]\[29\] registers\[31\]\[29\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__mux4_1
XFILLER_51_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35460_ clknet_leaf_231_CLK _03574_ VGND VGND VPWR VPWR registers\[14\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_16626_ registers\[32\]\[16\] registers\[33\]\[16\] registers\[34\]\[16\] registers\[35\]\[16\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15124_ sky130_fd_sc_hd__mux4_1
X_32672_ clknet_leaf_42_CLK _00786_ VGND VGND VPWR VPWR registers\[57\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34411_ clknet_leaf_401_CLK _02525_ VGND VGND VPWR VPWR registers\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_10_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_10_0_CLK sky130_fd_sc_hd__clkbuf_8
X_31623_ _14317_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__clkbuf_1
X_19345_ _06077_ _06080_ _05851_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35391_ clknet_leaf_297_CLK _03505_ VGND VGND VPWR VPWR registers\[15\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_16557_ _15034_ _15041_ _15050_ _15057_ VGND VGND VPWR VPWR _15058_ sky130_fd_sc_hd__or4_1
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34342_ clknet_leaf_448_CLK _02456_ VGND VGND VPWR VPWR registers\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31554_ _14281_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19276_ _05990_ _05997_ _06006_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__or4_4
XFILLER_203_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16488_ _14990_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18227_ _14600_ _04990_ _04991_ _14610_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__a22o_1
XFILLER_176_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30505_ _13729_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__clkbuf_1
X_34273_ clknet_leaf_41_CLK _02387_ VGND VGND VPWR VPWR registers\[32\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31485_ _09764_ registers\[6\]\[35\] _14239_ VGND VGND VPWR VPWR _14245_ sky130_fd_sc_hd__mux2_1
XFILLER_248_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_25_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_25_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_117_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36012_ clknet_leaf_374_CLK _04126_ VGND VGND VPWR VPWR registers\[63\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_33224_ clknet_leaf_211_CLK _01338_ VGND VGND VPWR VPWR registers\[4\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_30436_ _13637_ VGND VGND VPWR VPWR _13693_ sky130_fd_sc_hd__buf_4
X_18158_ registers\[44\]\[60\] registers\[45\]\[60\] registers\[46\]\[60\] registers\[47\]\[60\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__mux4_1
XFILLER_144_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17109_ _15487_ _15592_ _15593_ _15490_ VGND VGND VPWR VPWR _15594_ sky130_fd_sc_hd__a22o_1
X_33155_ clknet_leaf_270_CLK _01269_ VGND VGND VPWR VPWR registers\[50\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18089_ registers\[28\]\[57\] registers\[29\]\[57\] registers\[30\]\[57\] registers\[31\]\[57\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux4_1
X_30367_ _09693_ registers\[14\]\[17\] _13649_ VGND VGND VPWR VPWR _13657_ sky130_fd_sc_hd__mux2_1
X_20120_ registers\[28\]\[49\] registers\[29\]\[49\] registers\[30\]\[49\] registers\[31\]\[49\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32106_ clknet_leaf_483_CLK _00020_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33086_ clknet_leaf_267_CLK _01200_ VGND VGND VPWR VPWR registers\[51\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_30298_ registers\[15\]\[49\] _13037_ _13610_ VGND VGND VPWR VPWR _13620_ sky130_fd_sc_hd__mux2_1
XFILLER_131_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20051_ _06763_ _06766_ _06537_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__o21ba_1
X_32037_ clknet_leaf_450_CLK _00215_ VGND VGND VPWR VPWR registers\[62\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23810_ _09622_ registers\[29\]\[51\] _10072_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__mux2_1
XFILLER_26_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24790_ _09584_ registers\[54\]\[33\] _10620_ VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__mux2_1
X_33988_ clknet_leaf_252_CLK _02102_ VGND VGND VPWR VPWR registers\[37\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35727_ clknet_leaf_110_CLK _03841_ VGND VGND VPWR VPWR registers\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_20953_ _07281_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__clkbuf_4
X_23741_ _10037_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32939_ clknet_leaf_422_CLK _01053_ VGND VGND VPWR VPWR registers\[53\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26460_ _10775_ registers\[42\]\[21\] _11536_ VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__mux2_1
X_35658_ clknet_leaf_151_CLK _03772_ VGND VGND VPWR VPWR registers\[11\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_23672_ registers\[61\]\[51\] _09800_ _09998_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__mux2_1
X_20884_ _07333_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__clkbuf_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25411_ _10814_ registers\[50\]\[40\] _10981_ VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__mux2_1
X_22623_ registers\[4\]\[55\] registers\[5\]\[55\] registers\[6\]\[55\] registers\[7\]\[55\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__mux4_1
X_34609_ clknet_leaf_409_CLK _02723_ VGND VGND VPWR VPWR registers\[27\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_26391_ _11501_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35589_ clknet_leaf_227_CLK _03703_ VGND VGND VPWR VPWR registers\[12\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28130_ _11755_ registers\[30\]\[12\] _12446_ VGND VGND VPWR VPWR _12449_ sky130_fd_sc_hd__mux2_1
X_22554_ registers\[0\]\[53\] registers\[1\]\[53\] registers\[2\]\[53\] registers\[3\]\[53\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__mux4_1
X_25342_ _10945_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21505_ _08075_ _08179_ _08180_ _08078_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__a22o_1
X_28061_ _12412_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__clkbuf_1
X_22485_ registers\[8\]\[51\] registers\[9\]\[51\] registers\[10\]\[51\] registers\[11\]\[51\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__mux4_1
XFILLER_10_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25273_ _10908_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27012_ _11857_ registers\[3\]\[61\] _11729_ VGND VGND VPWR VPWR _11858_ sky130_fd_sc_hd__mux2_1
X_24224_ _09628_ registers\[58\]\[54\] _10288_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__mux2_1
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21436_ registers\[28\]\[21\] registers\[29\]\[21\] registers\[30\]\[21\] registers\[31\]\[21\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__mux4_1
XFILLER_181_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_17__f_CLK clknet_5_8_0_CLK VGND VGND VPWR VPWR clknet_6_17__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24155_ _09559_ registers\[58\]\[21\] _10255_ VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_190_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_190_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21367_ registers\[40\]\[20\] registers\[41\]\[20\] registers\[42\]\[20\] registers\[43\]\[20\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__mux4_1
XFILLER_174_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23106_ registers\[39\]\[6\] _09670_ _09658_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__mux2_1
X_20318_ _07022_ _07025_ _06855_ _06856_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__o211a_1
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24086_ _09626_ registers\[5\]\[53\] _10216_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__mux2_1
XFILLER_150_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28963_ registers\[24\]\[23\] _10353_ _12883_ VGND VGND VPWR VPWR _12887_ sky130_fd_sc_hd__mux2_1
X_21298_ registers\[44\]\[18\] registers\[45\]\[18\] registers\[46\]\[18\] registers\[47\]\[18\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__mux4_1
XFILLER_66_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23037_ _09621_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
X_27914_ registers\[32\]\[38\] _10384_ _12326_ VGND VGND VPWR VPWR _12335_ sky130_fd_sc_hd__mux2_1
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20249_ registers\[60\]\[53\] registers\[61\]\[53\] registers\[62\]\[53\] registers\[63\]\[53\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__mux4_1
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28894_ _12850_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__clkbuf_1
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27845_ registers\[32\]\[5\] _10315_ _12293_ VGND VGND VPWR VPWR _12299_ sky130_fd_sc_hd__mux2_1
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27776_ _12262_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__clkbuf_1
X_24988_ _10727_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__clkbuf_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29515_ _09823_ registers\[21\]\[62\] _13139_ VGND VGND VPWR VPWR _13208_ sky130_fd_sc_hd__mux2_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26727_ registers\[40\]\[19\] _10344_ _11669_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__mux2_1
XFILLER_205_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23939_ _09615_ registers\[60\]\[48\] _10133_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__mux2_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_710 _07301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_721 _07340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_732 _07352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29446_ _09751_ registers\[21\]\[29\] _13162_ VGND VGND VPWR VPWR _13172_ sky130_fd_sc_hd__mux2_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17460_ registers\[12\]\[39\] registers\[13\]\[39\] registers\[14\]\[39\] registers\[15\]\[39\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15935_ sky130_fd_sc_hd__mux4_1
XANTENNA_743 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26658_ _11642_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_754 _07385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_765 _07639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16411_ _14912_ _14915_ _14614_ VGND VGND VPWR VPWR _14916_ sky130_fd_sc_hd__o21ba_1
X_25609_ _11089_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_776 _08155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29377_ _13135_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_787 _08872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17391_ _15864_ _15867_ _15631_ VGND VGND VPWR VPWR _15868_ sky130_fd_sc_hd__o21ba_1
XFILLER_199_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_798 _08936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26589_ _10768_ registers\[41\]\[18\] _11597_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19130_ registers\[4\]\[21\] registers\[5\]\[21\] registers\[6\]\[21\] registers\[7\]\[21\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__mux4_1
X_16342_ registers\[40\]\[8\] registers\[41\]\[8\] registers\[42\]\[8\] registers\[43\]\[8\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14848_ sky130_fd_sc_hd__mux4_1
XFILLER_198_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28328_ registers\[2\]\[42\] _10393_ _12550_ VGND VGND VPWR VPWR _12553_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19061_ registers\[28\]\[19\] registers\[29\]\[19\] registers\[30\]\[19\] registers\[31\]\[19\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux4_1
XFILLER_12_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16273_ registers\[32\]\[6\] registers\[33\]\[6\] registers\[34\]\[6\] registers\[35\]\[6\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14781_ sky130_fd_sc_hd__mux4_1
X_28259_ _12516_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18012_ registers\[56\]\[55\] registers\[57\]\[55\] registers\[58\]\[55\] registers\[59\]\[55\]
+ _04751_ _04541_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__mux4_1
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31270_ _14131_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30221_ registers\[15\]\[12\] _12960_ _13577_ VGND VGND VPWR VPWR _13580_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_181_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_181_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30152_ _13543_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19963_ registers\[52\]\[45\] registers\[53\]\[45\] registers\[54\]\[45\] registers\[55\]\[45\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux4_1
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18914_ _05350_ _05660_ _05661_ _05353_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__a22o_1
XFILLER_84_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34960_ clknet_leaf_115_CLK _03074_ VGND VGND VPWR VPWR registers\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_30083_ _13507_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1120 _14573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19894_ registers\[48\]\[43\] registers\[49\]\[43\] registers\[50\]\[43\] registers\[51\]\[43\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__mux4_1
XTAP_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1131 _14607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1142 _14975_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1153 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33911_ clknet_leaf_336_CLK _02025_ VGND VGND VPWR VPWR registers\[38\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_18845_ _05069_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_1164 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34891_ clknet_leaf_143_CLK _03005_ VGND VGND VPWR VPWR registers\[23\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1175 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1186 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1197 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33842_ clknet_leaf_383_CLK _01956_ VGND VGND VPWR VPWR registers\[3\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_18776_ registers\[12\]\[11\] registers\[13\]\[11\] registers\[14\]\[11\] registers\[15\]\[11\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__mux4_1
X_15988_ _14492_ VGND VGND VPWR VPWR _14502_ sky130_fd_sc_hd__buf_12
XTAP_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17727_ _14573_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__clkbuf_4
XFILLER_76_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33773_ clknet_leaf_326_CLK _01887_ VGND VGND VPWR VPWR registers\[40\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_30985_ registers\[10\]\[54\] _13048_ _13977_ VGND VGND VPWR VPWR _13982_ sky130_fd_sc_hd__mux2_1
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35512_ clknet_leaf_320_CLK _03626_ VGND VGND VPWR VPWR registers\[13\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_32724_ clknet_leaf_65_CLK _00838_ VGND VGND VPWR VPWR registers\[56\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17658_ _04436_ _04439_ _15955_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16609_ registers\[8\]\[15\] registers\[9\]\[15\] registers\[10\]\[15\] registers\[11\]\[15\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15108_ sky130_fd_sc_hd__mux4_1
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32655_ clknet_leaf_75_CLK _00769_ VGND VGND VPWR VPWR registers\[57\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_35443_ clknet_leaf_354_CLK _03557_ VGND VGND VPWR VPWR registers\[14\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17589_ registers\[44\]\[43\] registers\[45\]\[43\] registers\[46\]\[43\] registers\[47\]\[43\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__mux4_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31606_ _14308_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__clkbuf_1
X_19328_ registers\[60\]\[27\] registers\[61\]\[27\] registers\[62\]\[27\] registers\[63\]\[27\]
+ _05962_ _05756_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__mux4_1
X_32586_ clknet_leaf_158_CLK _00700_ VGND VGND VPWR VPWR registers\[5\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35374_ clknet_leaf_393_CLK _03488_ VGND VGND VPWR VPWR registers\[15\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31537_ _09819_ registers\[6\]\[60\] _14205_ VGND VGND VPWR VPWR _14272_ sky130_fd_sc_hd__mux2_1
X_34325_ clknet_leaf_96_CLK _02439_ VGND VGND VPWR VPWR registers\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19259_ _05993_ _05996_ _05826_ _05827_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__o211a_1
XFILLER_149_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34256_ clknet_leaf_128_CLK _02370_ VGND VGND VPWR VPWR registers\[32\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_22270_ _08610_ _08922_ _08923_ _08613_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__a22o_1
XFILLER_129_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31468_ _09747_ registers\[6\]\[27\] _14228_ VGND VGND VPWR VPWR _14236_ sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33207_ clknet_leaf_313_CLK _01321_ VGND VGND VPWR VPWR registers\[4\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_21221_ _07737_ _07903_ _07904_ _07742_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__a22o_1
XFILLER_163_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30419_ _13684_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__clkbuf_1
X_34187_ clknet_leaf_158_CLK _02301_ VGND VGND VPWR VPWR registers\[34\]\[61\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_172_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_172_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31399_ _14199_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33138_ clknet_leaf_364_CLK _01252_ VGND VGND VPWR VPWR registers\[50\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_21152_ _07732_ _07836_ _07837_ _07735_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__a22o_1
XFILLER_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20103_ registers\[56\]\[49\] registers\[57\]\[49\] registers\[58\]\[49\] registers\[59\]\[49\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux4_1
X_25960_ _10814_ registers\[46\]\[40\] _11274_ VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__mux2_1
X_33069_ clknet_leaf_379_CLK _01183_ VGND VGND VPWR VPWR registers\[51\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_21083_ registers\[28\]\[11\] registers\[29\]\[11\] registers\[30\]\[11\] registers\[31\]\[11\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__mux4_1
XFILLER_59_814 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20034_ registers\[60\]\[47\] registers\[61\]\[47\] registers\[62\]\[47\] registers\[63\]\[47\]
+ _06648_ _06442_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__mux4_1
X_24911_ _10687_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25891_ _11238_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27630_ registers\[34\]\[31\] _10370_ _12184_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__mux2_1
X_24842_ _09636_ registers\[54\]\[58\] _10642_ VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__mux2_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27561_ _09867_ _10584_ VGND VGND VPWR VPWR _12148_ sky130_fd_sc_hd__or2_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24773_ _09567_ registers\[54\]\[25\] _10609_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__mux2_1
X_21985_ registers\[8\]\[37\] registers\[9\]\[37\] registers\[10\]\[37\] registers\[11\]\[37\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__mux4_1
X_29300_ _13095_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__clkbuf_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26512_ _10827_ registers\[42\]\[46\] _11558_ VGND VGND VPWR VPWR _11565_ sky130_fd_sc_hd__mux2_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23724_ _09535_ registers\[29\]\[10\] _10028_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__mux2_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ registers\[28\]\[7\] registers\[29\]\[7\] registers\[30\]\[7\] registers\[31\]\[7\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__mux4_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27492_ _12112_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29231_ net54 VGND VGND VPWR VPWR _13056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26443_ _10758_ registers\[42\]\[13\] _11525_ VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__mux2_1
XFILLER_187_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20867_ registers\[20\]\[5\] registers\[21\]\[5\] registers\[22\]\[5\] registers\[23\]\[5\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__mux4_1
XFILLER_169_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23655_ registers\[61\]\[43\] _09782_ _09987_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__mux2_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22606_ registers\[32\]\[55\] registers\[33\]\[55\] registers\[34\]\[55\] registers\[35\]\[55\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__mux4_1
XFILLER_224_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29162_ _13009_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26374_ _11492_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20798_ registers\[16\]\[3\] registers\[17\]\[3\] registers\[18\]\[3\] registers\[19\]\[3\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__mux4_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23586_ registers\[61\]\[10\] _09678_ _09954_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__mux2_1
X_28113_ _11738_ registers\[30\]\[4\] _12435_ VGND VGND VPWR VPWR _12440_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25325_ _10512_ _10935_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__nand2_8
XFILLER_122_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22537_ _09160_ _09167_ _09174_ _09183_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__or4_4
X_29093_ registers\[23\]\[13\] _12962_ _12956_ VGND VGND VPWR VPWR _12963_ sky130_fd_sc_hd__mux2_1
XFILLER_194_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28044_ _12403_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25256_ _10796_ registers\[51\]\[31\] _10898_ VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__mux2_1
X_22468_ _09108_ _09115_ _09116_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__o21ba_1
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24207_ _09611_ registers\[58\]\[46\] _10277_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_163_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_163_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21419_ registers\[56\]\[21\] registers\[57\]\[21\] registers\[58\]\[21\] registers\[59\]\[21\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__mux4_1
XFILLER_108_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25187_ _10862_ registers\[52\]\[63\] _10730_ VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__mux2_1
X_22399_ registers\[44\]\[49\] registers\[45\]\[49\] registers\[46\]\[49\] registers\[47\]\[49\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__mux4_1
XFILLER_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24138_ _09542_ registers\[58\]\[13\] _10244_ VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_1295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29995_ registers\[17\]\[33\] _13004_ _13457_ VGND VGND VPWR VPWR _13461_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16960_ _14502_ VGND VGND VPWR VPWR _15449_ sky130_fd_sc_hd__clkbuf_8
X_24069_ _09609_ registers\[5\]\[45\] _10205_ VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__mux2_1
X_28946_ registers\[24\]\[15\] _10336_ _12872_ VGND VGND VPWR VPWR _12878_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28877_ _12841_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__clkbuf_1
X_16891_ registers\[52\]\[23\] registers\[53\]\[23\] registers\[54\]\[23\] registers\[55\]\[23\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15382_ sky130_fd_sc_hd__mux4_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18630_ registers\[4\]\[7\] registers\[5\]\[7\] registers\[6\]\[7\] registers\[7\]\[7\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__mux4_1
X_27828_ _12289_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18561_ _05119_ _05317_ _05318_ _05131_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__a22o_1
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27759_ _12253_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17512_ _14581_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__clkbuf_4
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _05122_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__buf_4
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30770_ _09691_ registers\[11\]\[16\] _13862_ VGND VGND VPWR VPWR _13869_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_540 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_551 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_562 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17443_ _14520_ VGND VGND VPWR VPWR _15918_ sky130_fd_sc_hd__buf_4
X_29429_ _13163_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__clkbuf_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_573 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_584 _05067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_595 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32440_ clknet_leaf_429_CLK _00554_ VGND VGND VPWR VPWR registers\[29\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17374_ _14573_ VGND VGND VPWR VPWR _15851_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19113_ registers\[32\]\[21\] registers\[33\]\[21\] registers\[34\]\[21\] registers\[35\]\[21\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__mux4_1
XFILLER_159_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16325_ _14828_ _14831_ _14554_ _14556_ VGND VGND VPWR VPWR _14832_ sky130_fd_sc_hd__o211a_1
XFILLER_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32371_ clknet_leaf_357_CLK _00485_ VGND VGND VPWR VPWR registers\[61\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34110_ clknet_leaf_276_CLK _02224_ VGND VGND VPWR VPWR registers\[35\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31322_ _14159_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__clkbuf_1
X_19044_ registers\[56\]\[19\] registers\[57\]\[19\] registers\[58\]\[19\] registers\[59\]\[19\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__mux4_1
X_35090_ clknet_leaf_105_CLK _03204_ VGND VGND VPWR VPWR registers\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_16256_ registers\[8\]\[5\] registers\[9\]\[5\] registers\[10\]\[5\] registers\[11\]\[5\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14765_ sky130_fd_sc_hd__mux4_1
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34041_ clknet_leaf_337_CLK _02155_ VGND VGND VPWR VPWR registers\[36\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31253_ registers\[8\]\[53\] net49 _14119_ VGND VGND VPWR VPWR _14123_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_154_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_154_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16187_ _14694_ _14697_ _14554_ _14556_ VGND VGND VPWR VPWR _14698_ sky130_fd_sc_hd__o211a_1
XFILLER_154_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput205 net205 VGND VGND VPWR VPWR D2[56] sky130_fd_sc_hd__buf_2
XFILLER_245_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput216 net216 VGND VGND VPWR VPWR D2[8] sky130_fd_sc_hd__buf_2
X_30204_ registers\[15\]\[4\] _12943_ _13566_ VGND VGND VPWR VPWR _13571_ sky130_fd_sc_hd__mux2_1
Xoutput227 net227 VGND VGND VPWR VPWR D3[18] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR D3[28] sky130_fd_sc_hd__buf_2
XFILLER_177_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput249 net249 VGND VGND VPWR VPWR D3[38] sky130_fd_sc_hd__buf_2
X_31184_ registers\[8\]\[20\] net13 _14086_ VGND VGND VPWR VPWR _14087_ sky130_fd_sc_hd__mux2_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_63__f_CLK clknet_5_31_0_CLK VGND VGND VPWR VPWR clknet_6_63__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_30135_ _13534_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__clkbuf_1
X_19946_ registers\[28\]\[44\] registers\[29\]\[44\] registers\[30\]\[44\] registers\[31\]\[44\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__mux4_1
XFILLER_114_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35992_ clknet_leaf_58_CLK _04106_ VGND VGND VPWR VPWR registers\[63\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30066_ _13498_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__clkbuf_1
X_34943_ clknet_leaf_307_CLK _03057_ VGND VGND VPWR VPWR registers\[22\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_19877_ _06525_ _06596_ _06597_ _06528_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__a22o_1
XFILLER_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18828_ registers\[32\]\[13\] registers\[33\]\[13\] registers\[34\]\[13\] registers\[35\]\[13\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__mux4_1
X_34874_ clknet_leaf_309_CLK _02988_ VGND VGND VPWR VPWR registers\[23\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33825_ clknet_leaf_486_CLK _01939_ VGND VGND VPWR VPWR registers\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18759_ registers\[40\]\[11\] registers\[41\]\[11\] registers\[42\]\[11\] registers\[43\]\[11\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__mux4_1
X_21770_ _08126_ _08436_ _08437_ _08129_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__a22o_1
XFILLER_93_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30968_ registers\[10\]\[46\] _13031_ _13966_ VGND VGND VPWR VPWR _13973_ sky130_fd_sc_hd__mux2_1
X_33756_ clknet_leaf_28_CLK _01870_ VGND VGND VPWR VPWR registers\[40\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ registers\[0\]\[1\] registers\[1\]\[1\] registers\[2\]\[1\] registers\[3\]\[1\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__mux4_1
XFILLER_223_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32707_ clknet_leaf_270_CLK _00821_ VGND VGND VPWR VPWR registers\[57\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33687_ clknet_leaf_135_CLK _01801_ VGND VGND VPWR VPWR registers\[41\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_30899_ registers\[10\]\[13\] _12962_ _13933_ VGND VGND VPWR VPWR _13937_ sky130_fd_sc_hd__mux2_1
XFILLER_225_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20652_ registers\[0\]\[0\] registers\[1\]\[0\] registers\[2\]\[0\] registers\[3\]\[0\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__mux4_1
X_23440_ _09527_ registers\[19\]\[6\] _09870_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__mux2_1
X_35426_ clknet_leaf_467_CLK _03540_ VGND VGND VPWR VPWR registers\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_32638_ clknet_leaf_291_CLK _00752_ VGND VGND VPWR VPWR registers\[58\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23371_ registers\[39\]\[39\] _09773_ _09829_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__mux2_1
X_20583_ _07281_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__clkbuf_8
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32569_ clknet_leaf_315_CLK _00683_ VGND VGND VPWR VPWR registers\[5\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_35357_ clknet_leaf_480_CLK _03471_ VGND VGND VPWR VPWR registers\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_393_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_393_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25110_ _10810_ registers\[52\]\[38\] _10794_ VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__mux2_1
X_34308_ clknet_leaf_252_CLK _02422_ VGND VGND VPWR VPWR registers\[32\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_22322_ registers\[40\]\[47\] registers\[41\]\[47\] registers\[42\]\[47\] registers\[43\]\[47\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__mux4_1
X_26090_ _10810_ registers\[45\]\[38\] _11334_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35288_ clknet_leaf_8_CLK _03402_ VGND VGND VPWR VPWR registers\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22253_ registers\[32\]\[45\] registers\[33\]\[45\] registers\[34\]\[45\] registers\[35\]\[45\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__mux4_1
XFILLER_30_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25041_ net8 VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_145_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_145_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34239_ clknet_6_59__leaf_CLK _02353_ VGND VGND VPWR VPWR registers\[33\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21204_ registers\[52\]\[15\] registers\[53\]\[15\] registers\[54\]\[15\] registers\[55\]\[15\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__mux4_1
XFILLER_191_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22184_ _08817_ _08824_ _08831_ _08840_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__or4_4
XFILLER_172_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21135_ registers\[48\]\[13\] registers\[49\]\[13\] registers\[50\]\[13\] registers\[51\]\[13\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__mux4_1
X_28800_ _12789_ VGND VGND VPWR VPWR _12801_ sky130_fd_sc_hd__buf_4
X_29780_ _13347_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26992_ _11844_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28731_ _11816_ registers\[26\]\[41\] _12763_ VGND VGND VPWR VPWR _12765_ sky130_fd_sc_hd__mux2_1
XFILLER_87_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21066_ registers\[56\]\[11\] registers\[57\]\[11\] registers\[58\]\[11\] registers\[59\]\[11\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__mux4_1
XFILLER_115_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25943_ _10798_ registers\[46\]\[32\] _11263_ VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__mux2_1
XFILLER_87_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20017_ registers\[20\]\[46\] registers\[21\]\[46\] registers\[22\]\[46\] registers\[23\]\[46\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux4_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28662_ _12728_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25874_ _10585_ _11157_ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__nand2_8
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27613_ registers\[34\]\[23\] _10353_ _12173_ VGND VGND VPWR VPWR _12177_ sky130_fd_sc_hd__mux2_1
XFILLER_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24825_ _10586_ VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__clkbuf_8
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28593_ _12647_ VGND VGND VPWR VPWR _12692_ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27544_ _12139_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _09550_ registers\[54\]\[17\] _10598_ VGND VGND VPWR VPWR _10606_ sky130_fd_sc_hd__mux2_1
X_21968_ _08630_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__buf_6
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _09519_ registers\[29\]\[2\] _10017_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__mux2_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ registers\[56\]\[7\] registers\[57\]\[7\] registers\[58\]\[7\] registers\[59\]\[7\]
+ _07508_ _07317_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__mux4_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27475_ _12103_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_1
X_24687_ _10568_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21899_ registers\[40\]\[35\] registers\[41\]\[35\] registers\[42\]\[35\] registers\[43\]\[35\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__mux4_1
X_29214_ registers\[23\]\[52\] _13044_ _13040_ VGND VGND VPWR VPWR _13045_ sky130_fd_sc_hd__mux2_1
XFILLER_159_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26426_ _10741_ registers\[42\]\[5\] _11514_ VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__mux2_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ registers\[61\]\[35\] _09764_ _09976_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__mux2_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29145_ _12934_ VGND VGND VPWR VPWR _12998_ sky130_fd_sc_hd__buf_4
X_26357_ _11483_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__clkbuf_1
X_23569_ registers\[61\]\[2\] _09662_ _09943_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_384_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_384_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ registers\[36\]\[1\] registers\[37\]\[1\] registers\[38\]\[1\] registers\[39\]\[1\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14623_ sky130_fd_sc_hd__mux4_1
X_25308_ _10848_ registers\[51\]\[56\] _10920_ VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__mux2_1
XFILLER_156_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29076_ net63 VGND VGND VPWR VPWR _12951_ sky130_fd_sc_hd__clkbuf_4
X_17090_ _14520_ VGND VGND VPWR VPWR _15575_ sky130_fd_sc_hd__buf_4
X_26288_ _11447_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16041_ net70 VGND VGND VPWR VPWR _14555_ sky130_fd_sc_hd__buf_12
X_28027_ _12394_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_136_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_136_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_202_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25239_ _10779_ registers\[51\]\[23\] _10887_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19800_ _05133_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__buf_2
XFILLER_124_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17992_ _04486_ _04763_ _04764_ _04489_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__a22o_1
XFILLER_124_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29978_ registers\[17\]\[25\] _12987_ _13446_ VGND VGND VPWR VPWR _13452_ sky130_fd_sc_hd__mux2_1
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16943_ _15429_ _15432_ _15302_ VGND VGND VPWR VPWR _15433_ sky130_fd_sc_hd__o21ba_1
X_19731_ _06450_ _06455_ _06180_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__o21ba_1
X_28929_ registers\[24\]\[7\] _10319_ _12861_ VGND VGND VPWR VPWR _12869_ sky130_fd_sc_hd__mux2_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31940_ _09817_ registers\[49\]\[59\] _14474_ VGND VGND VPWR VPWR _14484_ sky130_fd_sc_hd__mux2_1
X_16874_ registers\[28\]\[22\] registers\[29\]\[22\] registers\[30\]\[22\] registers\[31\]\[22\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15366_ sky130_fd_sc_hd__mux4_1
X_19662_ _06182_ _06385_ _06388_ _06185_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__a22o_1
XFILLER_133_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18613_ registers\[44\]\[7\] registers\[45\]\[7\] registers\[46\]\[7\] registers\[47\]\[7\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ registers\[28\]\[34\] registers\[29\]\[34\] registers\[30\]\[34\] registers\[31\]\[34\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__mux4_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31871_ _09744_ registers\[49\]\[26\] _14441_ VGND VGND VPWR VPWR _14448_ sky130_fd_sc_hd__mux2_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33610_ clknet_leaf_161_CLK _01724_ VGND VGND VPWR VPWR registers\[43\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30822_ _13896_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__clkbuf_1
X_18544_ registers\[36\]\[5\] registers\[37\]\[5\] registers\[38\]\[5\] registers\[39\]\[5\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__mux4_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34590_ clknet_leaf_4_CLK _02704_ VGND VGND VPWR VPWR registers\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18475_ registers\[32\]\[3\] registers\[33\]\[3\] registers\[34\]\[3\] registers\[35\]\[3\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__mux4_1
X_33541_ clknet_leaf_256_CLK _01655_ VGND VGND VPWR VPWR registers\[44\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_30753_ _09674_ registers\[11\]\[8\] _13851_ VGND VGND VPWR VPWR _13860_ sky130_fd_sc_hd__mux2_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_370 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_381 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17426_ registers\[12\]\[38\] registers\[13\]\[38\] registers\[14\]\[38\] registers\[15\]\[38\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15902_ sky130_fd_sc_hd__mux4_1
X_33472_ clknet_leaf_256_CLK _01586_ VGND VGND VPWR VPWR registers\[45\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30684_ _13823_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35211_ clknet_leaf_149_CLK _03325_ VGND VGND VPWR VPWR registers\[18\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32423_ clknet_leaf_456_CLK _00537_ VGND VGND VPWR VPWR registers\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17357_ _15829_ _15834_ _15631_ VGND VGND VPWR VPWR _15835_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36191_ clknet_leaf_29_CLK _00072_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_375_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_375_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16308_ _14786_ _14795_ _14806_ _14815_ VGND VGND VPWR VPWR _14816_ sky130_fd_sc_hd__or4_4
X_35142_ clknet_leaf_217_CLK _03256_ VGND VGND VPWR VPWR registers\[1\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_32354_ clknet_leaf_444_CLK _00468_ VGND VGND VPWR VPWR registers\[61\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17288_ _14562_ VGND VGND VPWR VPWR _15768_ sky130_fd_sc_hd__buf_6
XFILLER_88_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19027_ registers\[16\]\[18\] registers\[17\]\[18\] registers\[18\]\[18\] registers\[19\]\[18\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__mux4_1
X_31305_ _14150_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__clkbuf_1
X_35073_ clknet_leaf_202_CLK _03187_ VGND VGND VPWR VPWR registers\[20\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_16239_ _14748_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_127_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_127_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32285_ clknet_leaf_5_CLK _00399_ VGND VGND VPWR VPWR registers\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34024_ clknet_leaf_435_CLK _02138_ VGND VGND VPWR VPWR registers\[36\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31236_ registers\[8\]\[45\] net40 _14108_ VGND VGND VPWR VPWR _14114_ sky130_fd_sc_hd__mux2_1
XFILLER_6_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31167_ registers\[8\]\[12\] net4 _14075_ VGND VGND VPWR VPWR _14078_ sky130_fd_sc_hd__mux2_1
XFILLER_88_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30118_ _13525_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__clkbuf_1
X_19929_ _05090_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__buf_6
XFILLER_69_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35975_ clknet_leaf_210_CLK _04089_ VGND VGND VPWR VPWR registers\[6\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_31098_ _14041_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30049_ registers\[17\]\[59\] _13058_ _13479_ VGND VGND VPWR VPWR _13489_ sky130_fd_sc_hd__mux2_1
X_34926_ clknet_leaf_394_CLK _03040_ VGND VGND VPWR VPWR registers\[22\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_22940_ _09555_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22871_ _07355_ _09505_ _09506_ _07367_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__a22o_1
X_34857_ clknet_leaf_454_CLK _02971_ VGND VGND VPWR VPWR registers\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24610_ _10528_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33808_ clknet_leaf_111_CLK _01922_ VGND VGND VPWR VPWR registers\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_21822_ registers\[24\]\[32\] registers\[25\]\[32\] registers\[26\]\[32\] registers\[27\]\[32\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__mux4_1
XFILLER_225_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25590_ _11077_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34788_ clknet_leaf_446_CLK _02902_ VGND VGND VPWR VPWR registers\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24541_ _10490_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33739_ clknet_leaf_156_CLK _01853_ VGND VGND VPWR VPWR registers\[41\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_21753_ _08418_ _08419_ _08420_ _08421_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__a22o_1
XFILLER_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20704_ registers\[40\]\[1\] registers\[41\]\[1\] registers\[42\]\[1\] registers\[43\]\[1\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__mux4_1
X_27260_ _11832_ registers\[37\]\[49\] _11980_ VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__mux2_1
X_24472_ _10454_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21684_ _08080_ _08353_ _08354_ _08085_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__a22o_1
XFILLER_221_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26211_ _10796_ registers\[44\]\[31\] _11405_ VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__mux2_1
X_23423_ _09651_ _09650_ _09649_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__nor3b_4
X_35409_ clknet_leaf_107_CLK _03523_ VGND VGND VPWR VPWR registers\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20635_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_366_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_366_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27191_ _11763_ registers\[37\]\[16\] _11947_ VGND VGND VPWR VPWR _11954_ sky130_fd_sc_hd__mux2_1
XFILLER_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26142_ _10862_ registers\[45\]\[63\] _11300_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__mux2_1
X_20566_ registers\[24\]\[63\] registers\[25\]\[63\] registers\[26\]\[63\] registers\[27\]\[63\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__mux4_1
X_23354_ _09830_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22305_ _07295_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_118_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_118_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26073_ _11300_ VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__buf_4
X_20497_ _05149_ _07197_ _07198_ _05159_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__a22o_1
X_23285_ _09785_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29901_ _13411_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__clkbuf_1
X_25024_ _10751_ registers\[52\]\[10\] _10752_ VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22236_ _08610_ _08889_ _08890_ _08613_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__a22o_1
XFILLER_69_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22167_ _08820_ _08823_ _08748_ _08749_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__o211a_1
X_29832_ _13352_ VGND VGND VPWR VPWR _13375_ sky130_fd_sc_hd__buf_4
XTAP_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1708 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1719 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21118_ _07732_ _07803_ _07804_ _07735_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__a22o_1
XTAP_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29763_ registers\[1\]\[51\] _13042_ _13337_ VGND VGND VPWR VPWR _13339_ sky130_fd_sc_hd__mux2_1
X_26975_ _11832_ registers\[3\]\[49\] _11814_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__mux2_1
X_22098_ registers\[4\]\[40\] registers\[5\]\[40\] registers\[6\]\[40\] registers\[7\]\[40\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__mux4_1
XTAP_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25926_ _10781_ registers\[46\]\[24\] _11252_ VGND VGND VPWR VPWR _11257_ sky130_fd_sc_hd__mux2_1
X_28714_ _11799_ registers\[26\]\[33\] _12752_ VGND VGND VPWR VPWR _12756_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21049_ registers\[28\]\[10\] registers\[29\]\[10\] registers\[30\]\[10\] registers\[31\]\[10\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__mux4_1
X_29694_ _13302_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28645_ _11728_ registers\[26\]\[0\] _12719_ VGND VGND VPWR VPWR _12720_ sky130_fd_sc_hd__mux2_1
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25857_ _11220_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24808_ _10633_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
X_28576_ _12683_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__clkbuf_1
X_16590_ _15086_ _15089_ _14959_ VGND VGND VPWR VPWR _15090_ sky130_fd_sc_hd__o21ba_1
X_25788_ _11184_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27527_ _12130_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__clkbuf_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24739_ _09533_ registers\[54\]\[9\] _10587_ VGND VGND VPWR VPWR _10597_ sky130_fd_sc_hd__mux2_1
XFILLER_131_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ registers\[0\]\[63\] registers\[1\]\[63\] registers\[2\]\[63\] registers\[3\]\[63\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__mux4_1
XFILLER_230_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27458_ _12094_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ registers\[60\]\[32\] registers\[61\]\[32\] registers\[62\]\[32\] registers\[63\]\[32\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15693_ sky130_fd_sc_hd__mux4_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26409_ _11510_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__clkbuf_1
X_18191_ _04953_ _04956_ _14524_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__o21ba_1
XFILLER_202_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27389_ registers\[36\]\[46\] _10401_ _12051_ VGND VGND VPWR VPWR _12058_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_357_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_357_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17142_ registers\[0\]\[30\] registers\[1\]\[30\] registers\[2\]\[30\] registers\[3\]\[30\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15626_ sky130_fd_sc_hd__mux4_1
X_29128_ _12986_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29059_ registers\[23\]\[2\] _12939_ _12935_ VGND VGND VPWR VPWR _12940_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_109_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_109_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17073_ registers\[12\]\[28\] registers\[13\]\[28\] registers\[14\]\[28\] registers\[15\]\[28\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15559_ sky130_fd_sc_hd__mux4_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16024_ _14528_ _14533_ _14536_ _14537_ VGND VGND VPWR VPWR _14538_ sky130_fd_sc_hd__a22o_1
X_32070_ clknet_leaf_194_CLK _00248_ VGND VGND VPWR VPWR registers\[62\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31021_ registers\[0\]\[7\] _12949_ _13993_ VGND VGND VPWR VPWR _14001_ sky130_fd_sc_hd__mux2_1
XFILLER_156_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17975_ registers\[36\]\[54\] registers\[37\]\[54\] registers\[38\]\[54\] registers\[39\]\[54\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux4_1
XFILLER_112_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19714_ _05049_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__clkbuf_4
X_35760_ clknet_leaf_377_CLK _03874_ VGND VGND VPWR VPWR registers\[0\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_16926_ _15206_ _15414_ _15415_ _15210_ VGND VGND VPWR VPWR _15416_ sky130_fd_sc_hd__a22o_1
X_32972_ clknet_leaf_142_CLK _01086_ VGND VGND VPWR VPWR registers\[53\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34711_ clknet_leaf_94_CLK _02825_ VGND VGND VPWR VPWR registers\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_31923_ _14475_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_1
X_19645_ _06098_ _06368_ _06371_ _06102_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__a22o_1
X_35691_ clknet_leaf_399_CLK _03805_ VGND VGND VPWR VPWR registers\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16857_ _15198_ _15347_ _15348_ _15204_ VGND VGND VPWR VPWR _15349_ sky130_fd_sc_hd__a22o_1
XFILLER_168_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34642_ clknet_leaf_95_CLK _02756_ VGND VGND VPWR VPWR registers\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16788_ _14564_ VGND VGND VPWR VPWR _15282_ sky130_fd_sc_hd__clkbuf_4
X_31854_ _09695_ registers\[49\]\[18\] _14430_ VGND VGND VPWR VPWR _14439_ sky130_fd_sc_hd__mux2_1
X_19576_ _05090_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__buf_6
XFILLER_20_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18527_ _05119_ _05284_ _05285_ _05131_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__a22o_1
X_30805_ _13887_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34573_ clknet_leaf_140_CLK _02687_ VGND VGND VPWR VPWR registers\[28\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_31785_ _14402_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33524_ clknet_leaf_346_CLK _01638_ VGND VGND VPWR VPWR registers\[44\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_18458_ _05107_ _05217_ _05218_ _05117_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__a22o_1
X_30736_ _13850_ VGND VGND VPWR VPWR _13851_ sky130_fd_sc_hd__buf_4
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17409_ _14531_ VGND VGND VPWR VPWR _15885_ sky130_fd_sc_hd__buf_4
X_18389_ _05080_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__buf_12
X_30667_ registers\[12\]\[31\] _13000_ _13813_ VGND VGND VPWR VPWR _13815_ sky130_fd_sc_hd__mux2_1
X_33455_ clknet_leaf_363_CLK _01569_ VGND VGND VPWR VPWR registers\[45\]\[33\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_348_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_348_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20420_ registers\[20\]\[58\] registers\[21\]\[58\] registers\[22\]\[58\] registers\[23\]\[58\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__mux4_1
XFILLER_53_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32406_ clknet_leaf_88_CLK _00520_ VGND VGND VPWR VPWR registers\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_36174_ clknet_leaf_92_CLK _00064_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_1
X_30598_ _09825_ registers\[13\]\[63\] _13708_ VGND VGND VPWR VPWR _13778_ sky130_fd_sc_hd__mux2_1
X_33386_ clknet_leaf_429_CLK _01500_ VGND VGND VPWR VPWR registers\[46\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20351_ _05040_ _07056_ _07057_ _05050_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__a22o_1
X_35125_ clknet_leaf_383_CLK _03239_ VGND VGND VPWR VPWR registers\[1\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_32337_ clknet_leaf_180_CLK _00451_ VGND VGND VPWR VPWR registers\[61\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23070_ _09643_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
X_32268_ clknet_leaf_168_CLK _00382_ VGND VGND VPWR VPWR registers\[39\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_20282_ _05090_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__buf_6
X_35056_ clknet_leaf_389_CLK _03170_ VGND VGND VPWR VPWR registers\[20\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22021_ _08677_ _08679_ _08680_ _08681_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__a22o_1
XTAP_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34007_ clknet_leaf_119_CLK _02121_ VGND VGND VPWR VPWR registers\[36\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_31219_ registers\[8\]\[37\] net31 _14097_ VGND VGND VPWR VPWR _14105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32199_ clknet_leaf_391_CLK _00313_ VGND VGND VPWR VPWR registers\[9\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26760_ _11696_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__clkbuf_1
X_23972_ _09651_ _09649_ _09650_ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__nor3_4
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35958_ clknet_leaf_319_CLK _04072_ VGND VGND VPWR VPWR registers\[6\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_25711_ registers\[48\]\[51\] _10412_ _11141_ VGND VGND VPWR VPWR _11143_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34909_ clknet_leaf_491_CLK _03023_ VGND VGND VPWR VPWR registers\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_22923_ net6 VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__buf_4
X_26691_ _11660_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__clkbuf_1
X_35889_ clknet_leaf_374_CLK _04003_ VGND VGND VPWR VPWR registers\[7\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28430_ _12606_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25642_ _11106_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22854_ _07372_ _09488_ _09489_ _07382_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__a22o_1
XFILLER_56_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28361_ registers\[2\]\[58\] _10426_ _12561_ VGND VGND VPWR VPWR _12570_ sky130_fd_sc_hd__mux2_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21805_ _07301_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__clkbuf_4
X_25573_ registers\[4\]\[51\] _10412_ _11067_ VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__mux2_1
XFILLER_71_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22785_ registers\[40\]\[61\] registers\[41\]\[61\] registers\[42\]\[61\] registers\[43\]\[61\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__mux4_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27312_ _12017_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__clkbuf_1
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24524_ _10481_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28292_ registers\[2\]\[25\] _10357_ _12528_ VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__mux2_1
XFILLER_40_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21736_ _07338_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__clkbuf_4
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27243_ _11981_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24455_ _10445_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_339_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_339_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21667_ _07301_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23406_ _09857_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
X_27174_ _11746_ registers\[37\]\[8\] _11936_ VGND VGND VPWR VPWR _11945_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20618_ _07316_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__buf_4
XFILLER_123_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24386_ registers\[57\]\[45\] _10399_ _10389_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21598_ _08267_ _08268_ _08269_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__a22o_1
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26125_ _11361_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23337_ registers\[9\]\[60\] _09819_ _09708_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20549_ registers\[36\]\[63\] registers\[37\]\[63\] registers\[38\]\[63\] registers\[39\]\[63\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__mux4_1
XFILLER_197_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26056_ _11325_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
X_23268_ registers\[9\]\[39\] _09773_ _09754_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__mux2_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25007_ net56 VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__buf_4
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22219_ registers\[32\]\[44\] registers\[33\]\[44\] registers\[34\]\[44\] registers\[35\]\[44\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__mux4_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23199_ net16 VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__clkbuf_4
XTAP_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1505 _07382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1516 _08668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1527 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29815_ _13366_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1538 _09780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1549 _10749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17760_ _04535_ _04538_ _15955_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__o21ba_1
X_29746_ registers\[1\]\[43\] _13025_ _13326_ VGND VGND VPWR VPWR _13330_ sky130_fd_sc_hd__mux2_1
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26958_ _11821_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_873 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16711_ _14543_ VGND VGND VPWR VPWR _15207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_248_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17691_ registers\[56\]\[46\] registers\[57\]\[46\] registers\[58\]\[46\] registers\[59\]\[46\]
+ _04408_ _15885_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__mux4_1
XFILLER_101_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25909_ _10764_ registers\[46\]\[16\] _11241_ VGND VGND VPWR VPWR _11248_ sky130_fd_sc_hd__mux2_1
XFILLER_235_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26889_ _11774_ registers\[3\]\[21\] _11772_ VGND VGND VPWR VPWR _11775_ sky130_fd_sc_hd__mux2_1
X_29677_ registers\[1\]\[10\] _12955_ _13293_ VGND VGND VPWR VPWR _13294_ sky130_fd_sc_hd__mux2_1
XFILLER_207_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19430_ registers\[56\]\[30\] registers\[57\]\[30\] registers\[58\]\[30\] registers\[59\]\[30\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__mux4_1
X_16642_ registers\[8\]\[16\] registers\[9\]\[16\] registers\[10\]\[16\] registers\[11\]\[16\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15140_ sky130_fd_sc_hd__mux4_1
X_28628_ _12710_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19361_ _05049_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__clkbuf_8
X_16573_ _14863_ _15071_ _15072_ _14867_ VGND VGND VPWR VPWR _15073_ sky130_fd_sc_hd__a22o_1
X_28559_ _12674_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__clkbuf_1
X_18312_ _05056_ _05072_ _05074_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__o21ba_1
XFILLER_206_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31570_ registers\[63\]\[11\] net3 _14288_ VGND VGND VPWR VPWR _14290_ sky130_fd_sc_hd__mux2_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _05755_ _06025_ _06028_ _05759_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__a22o_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _04986_ _04993_ _05000_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__or4_4
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30521_ _09744_ registers\[13\]\[26\] _13731_ VGND VGND VPWR VPWR _13738_ sky130_fd_sc_hd__mux2_1
XFILLER_175_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18174_ _14511_ _04939_ _04940_ _14517_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__a22o_1
X_30452_ _13701_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33240_ clknet_leaf_51_CLK _01354_ VGND VGND VPWR VPWR registers\[48\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17125_ registers\[44\]\[30\] registers\[45\]\[30\] registers\[46\]\[30\] registers\[47\]\[30\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15609_ sky130_fd_sc_hd__mux4_2
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33171_ clknet_leaf_78_CLK _01285_ VGND VGND VPWR VPWR registers\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30383_ _13665_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32122_ clknet_leaf_393_CLK _00038_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17056_ _14531_ VGND VGND VPWR VPWR _15542_ sky130_fd_sc_hd__buf_6
X_16007_ _14520_ VGND VGND VPWR VPWR _14521_ sky130_fd_sc_hd__buf_4
X_32053_ clknet_leaf_325_CLK _00231_ VGND VGND VPWR VPWR registers\[62\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31004_ _13991_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__clkbuf_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35812_ clknet_leaf_465_CLK _03926_ VGND VGND VPWR VPWR registers\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ registers\[12\]\[53\] registers\[13\]\[53\] registers\[14\]\[53\] registers\[15\]\[53\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__mux4_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35743_ clknet_leaf_486_CLK _03857_ VGND VGND VPWR VPWR registers\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16909_ _15396_ _15399_ _15302_ VGND VGND VPWR VPWR _15400_ sky130_fd_sc_hd__o21ba_1
X_32955_ clknet_leaf_287_CLK _01069_ VGND VGND VPWR VPWR registers\[53\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_17889_ registers\[4\]\[51\] registers\[5\]\[51\] registers\[6\]\[51\] registers\[7\]\[51\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__mux4_1
XFILLER_96_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31906_ _14466_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__clkbuf_1
X_19628_ _06352_ _06355_ _06194_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__o21ba_1
X_35674_ clknet_leaf_15_CLK _03788_ VGND VGND VPWR VPWR registers\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_32886_ clknet_leaf_326_CLK _01000_ VGND VGND VPWR VPWR registers\[54\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34625_ clknet_leaf_222_CLK _02739_ VGND VGND VPWR VPWR registers\[27\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19559_ registers\[28\]\[33\] registers\[29\]\[33\] registers\[30\]\[33\] registers\[31\]\[33\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__mux4_1
X_31837_ _14418_ VGND VGND VPWR VPWR _14430_ sky130_fd_sc_hd__buf_4
XFILLER_202_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22570_ _09215_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34556_ clknet_leaf_187_CLK _02670_ VGND VGND VPWR VPWR registers\[28\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_31768_ registers\[59\]\[41\] net36 _14392_ VGND VGND VPWR VPWR _14394_ sky130_fd_sc_hd__mux2_1
XFILLER_222_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33507_ clknet_leaf_59_CLK _01621_ VGND VGND VPWR VPWR registers\[44\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_21521_ registers\[48\]\[24\] registers\[49\]\[24\] registers\[50\]\[24\] registers\[51\]\[24\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__mux4_1
X_30719_ registers\[12\]\[56\] _13052_ _13835_ VGND VGND VPWR VPWR _13842_ sky130_fd_sc_hd__mux2_1
XFILLER_178_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34487_ clknet_leaf_314_CLK _02601_ VGND VGND VPWR VPWR registers\[2\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31699_ _14357_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36226_ clknet_leaf_121_CLK _00111_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dfxtp_1
X_24240_ _09644_ registers\[58\]\[62\] _10232_ VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__mux2_1
XFILLER_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21452_ _07301_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__buf_4
X_33438_ clknet_leaf_26_CLK _01552_ VGND VGND VPWR VPWR registers\[45\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_20403_ registers\[48\]\[58\] registers\[49\]\[58\] registers\[50\]\[58\] registers\[51\]\[58\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__mux4_1
X_36157_ clknet_leaf_290_CLK _04271_ VGND VGND VPWR VPWR registers\[49\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21383_ _07338_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__clkbuf_4
X_24171_ _09575_ registers\[58\]\[29\] _10255_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__mux2_1
X_33369_ clknet_leaf_29_CLK _01483_ VGND VGND VPWR VPWR registers\[46\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23122_ registers\[39\]\[11\] _09681_ _09679_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__mux2_1
X_35108_ clknet_leaf_465_CLK _03222_ VGND VGND VPWR VPWR registers\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_20334_ _07041_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__buf_4
XFILLER_134_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36088_ clknet_leaf_334_CLK _04202_ VGND VGND VPWR VPWR registers\[59\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20265_ registers\[28\]\[53\] registers\[29\]\[53\] registers\[30\]\[53\] registers\[31\]\[53\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__mux4_1
XFILLER_190_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23053_ net52 VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__clkbuf_8
X_27930_ _12343_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__clkbuf_1
X_35039_ clknet_leaf_489_CLK _03153_ VGND VGND VPWR VPWR registers\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22004_ registers\[44\]\[38\] registers\[45\]\[38\] registers\[46\]\[38\] registers\[47\]\[38\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__mux4_1
XFILLER_248_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27861_ _12307_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20196_ registers\[20\]\[51\] registers\[21\]\[51\] registers\[22\]\[51\] registers\[23\]\[51\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux4_1
XTAP_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29600_ registers\[20\]\[38\] _13014_ _13244_ VGND VGND VPWR VPWR _13253_ sky130_fd_sc_hd__mux2_1
X_26812_ _11723_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_1
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27792_ registers\[33\]\[44\] _10397_ _12266_ VGND VGND VPWR VPWR _12271_ sky130_fd_sc_hd__mux2_1
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29531_ registers\[20\]\[5\] _12945_ _13211_ VGND VGND VPWR VPWR _13217_ sky130_fd_sc_hd__mux2_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26743_ _11687_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__clkbuf_1
X_23955_ _10150_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22906_ _09532_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29462_ _13180_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__clkbuf_1
X_26674_ _11650_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_903 _09660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23886_ _10114_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_914 _09708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_925 _09815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25625_ registers\[48\]\[10\] _10325_ _11097_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__mux2_1
XFILLER_112_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28413_ _12597_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_936 _10160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22837_ registers\[16\]\[62\] registers\[17\]\[62\] registers\[18\]\[62\] registers\[19\]\[62\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__mux4_1
X_29393_ _13144_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_947 _10391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_958 _10796_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_969 _10936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28344_ _12505_ VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__buf_4
XFILLER_164_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25556_ registers\[4\]\[43\] _10395_ _11056_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__mux2_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22768_ _09403_ _09406_ _07338_ _07340_ VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__o211a_1
XFILLER_38_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24507_ _10472_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28275_ registers\[2\]\[17\] _10340_ _12517_ VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__mux2_1
X_21719_ _08388_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25487_ registers\[4\]\[10\] _10325_ _11023_ VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__mux2_1
X_22699_ registers\[36\]\[58\] registers\[37\]\[58\] registers\[38\]\[58\] registers\[39\]\[58\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__mux4_1
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27226_ _11972_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__clkbuf_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24438_ registers\[57\]\[62\] _10434_ net283 VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__mux2_1
XFILLER_138_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27157_ _11935_ VGND VGND VPWR VPWR _11936_ sky130_fd_sc_hd__buf_4
X_24369_ net35 VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__clkbuf_4
X_26108_ _11352_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27088_ _11795_ registers\[38\]\[31\] _11898_ VGND VGND VPWR VPWR _11900_ sky130_fd_sc_hd__mux2_1
XFILLER_180_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26039_ _11316_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
X_18930_ _05547_ _05675_ _05676_ _05550_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__a22o_1
XFILLER_238_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_40_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1302 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1313 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18861_ _05540_ _05608_ _05609_ _05545_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__a22o_1
XTAP_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1324 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1335 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1346 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17812_ _04481_ _04588_ _04589_ _04484_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__a22o_1
XFILLER_121_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1357 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1368 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18792_ registers\[40\]\[12\] registers\[41\]\[12\] registers\[42\]\[12\] registers\[43\]\[12\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__mux4_1
XFILLER_239_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1379 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _04486_ _04521_ _04522_ _04489_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__a22o_1
X_29729_ registers\[1\]\[35\] _13008_ _13315_ VGND VGND VPWR VPWR _13321_ sky130_fd_sc_hd__mux2_1
XFILLER_36_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32740_ clknet_leaf_441_CLK _00854_ VGND VGND VPWR VPWR registers\[56\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_17674_ _04452_ _04455_ _15974_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__o21ba_1
XFILLER_75_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19413_ _05839_ _06145_ _06146_ _05842_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__a22o_1
XFILLER_78_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16625_ registers\[40\]\[16\] registers\[41\]\[16\] registers\[42\]\[16\] registers\[43\]\[16\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15123_ sky130_fd_sc_hd__mux4_1
X_32671_ clknet_leaf_38_CLK _00785_ VGND VGND VPWR VPWR registers\[57\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34410_ clknet_leaf_404_CLK _02524_ VGND VGND VPWR VPWR registers\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19344_ _05844_ _06078_ _06079_ _05849_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__a22o_1
X_31622_ registers\[63\]\[36\] net30 _14310_ VGND VGND VPWR VPWR _14317_ sky130_fd_sc_hd__mux2_1
X_16556_ _15053_ _15056_ _14959_ VGND VGND VPWR VPWR _15057_ sky130_fd_sc_hd__o21ba_1
X_35390_ clknet_leaf_197_CLK _03504_ VGND VGND VPWR VPWR registers\[15\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34341_ clknet_leaf_464_CLK _02455_ VGND VGND VPWR VPWR registers\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_31553_ registers\[63\]\[3\] net34 _14277_ VGND VGND VPWR VPWR _14281_ sky130_fd_sc_hd__mux2_1
X_19275_ _06009_ _06012_ _05851_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__o21ba_1
X_16487_ _14968_ _14975_ _14982_ _14989_ VGND VGND VPWR VPWR _14990_ sky130_fd_sc_hd__or4_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18226_ registers\[52\]\[62\] registers\[53\]\[62\] registers\[54\]\[62\] registers\[55\]\[62\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__mux4_1
X_30504_ _09695_ registers\[13\]\[18\] _13720_ VGND VGND VPWR VPWR _13729_ sky130_fd_sc_hd__mux2_1
X_31484_ _14244_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__clkbuf_1
X_34272_ clknet_leaf_17_CLK _02386_ VGND VGND VPWR VPWR registers\[32\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36011_ clknet_leaf_422_CLK _04125_ VGND VGND VPWR VPWR registers\[63\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_33223_ clknet_leaf_210_CLK _01337_ VGND VGND VPWR VPWR registers\[4\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_30435_ _13692_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__clkbuf_1
X_18157_ _04676_ _04922_ _04923_ _04681_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__a22o_1
XFILLER_157_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17108_ registers\[4\]\[29\] registers\[5\]\[29\] registers\[6\]\[29\] registers\[7\]\[29\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15593_ sky130_fd_sc_hd__mux4_1
X_18088_ _04632_ _04856_ _04857_ _04635_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a22o_1
X_33154_ clknet_leaf_263_CLK _01268_ VGND VGND VPWR VPWR registers\[50\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30366_ _13656_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32105_ clknet_leaf_483_CLK _00019_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dfxtp_1
X_17039_ registers\[24\]\[27\] registers\[25\]\[27\] registers\[26\]\[27\] registers\[27\]\[27\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15526_ sky130_fd_sc_hd__mux4_1
X_33085_ clknet_leaf_268_CLK _01199_ VGND VGND VPWR VPWR registers\[51\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_30297_ _13619_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_31_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_31_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20050_ _06530_ _06764_ _06765_ _06535_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a22o_1
X_32036_ clknet_leaf_446_CLK _00214_ VGND VGND VPWR VPWR registers\[62\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33987_ clknet_leaf_252_CLK _02101_ VGND VGND VPWR VPWR registers\[37\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35726_ clknet_leaf_110_CLK _03840_ VGND VGND VPWR VPWR registers\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_23740_ _09552_ registers\[29\]\[18\] _10028_ VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__mux2_1
XFILLER_27_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _07278_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__buf_4
X_32938_ clknet_leaf_407_CLK _01052_ VGND VGND VPWR VPWR registers\[53\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35657_ clknet_leaf_155_CLK _03771_ VGND VGND VPWR VPWR registers\[11\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23671_ _09999_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_98_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_98_CLK sky130_fd_sc_hd__clkbuf_16
X_20883_ _07331_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__buf_4
X_32869_ clknet_leaf_438_CLK _00983_ VGND VGND VPWR VPWR registers\[54\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25410_ _10936_ VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__buf_4
X_22622_ registers\[12\]\[55\] registers\[13\]\[55\] registers\[14\]\[55\] registers\[15\]\[55\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__mux4_1
XFILLER_35_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34608_ clknet_leaf_411_CLK _02722_ VGND VGND VPWR VPWR registers\[27\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_26390_ _10840_ registers\[43\]\[52\] _11498_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__mux2_1
X_35588_ clknet_leaf_231_CLK _03702_ VGND VGND VPWR VPWR registers\[12\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25341_ _10745_ registers\[50\]\[7\] _10937_ VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__mux2_1
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22553_ registers\[8\]\[53\] registers\[9\]\[53\] registers\[10\]\[53\] registers\[11\]\[53\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__mux4_1
X_34539_ clknet_leaf_401_CLK _02653_ VGND VGND VPWR VPWR registers\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28060_ _11820_ registers\[31\]\[43\] _12408_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__mux2_1
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21504_ registers\[16\]\[23\] registers\[17\]\[23\] registers\[18\]\[23\] registers\[19\]\[23\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__mux4_1
X_25272_ _10812_ registers\[51\]\[39\] _10898_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__mux2_1
X_22484_ _09128_ _09131_ _09091_ _09092_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__o211a_1
XFILLER_210_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27011_ net58 VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__buf_2
XFILLER_194_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36209_ clknet_leaf_115_CLK _00092_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dfxtp_1
X_24223_ _10292_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21435_ _08075_ _08111_ _08112_ _08078_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__a22o_1
XFILLER_198_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24154_ _10256_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
X_21366_ _08045_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23105_ net61 VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__buf_4
X_20317_ _06784_ _07023_ _07024_ _06788_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__a22o_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24085_ _10219_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28962_ _12886_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_22_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_22_CLK sky130_fd_sc_hd__clkbuf_16
X_21297_ _07776_ _07976_ _07977_ _07781_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__a22o_1
X_23036_ _09619_ registers\[62\]\[50\] _09620_ VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__mux2_1
X_27913_ _12334_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20248_ _06776_ _06956_ _06957_ _06782_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__a22o_1
X_28893_ _11843_ registers\[25\]\[54\] _12845_ VGND VGND VPWR VPWR _12850_ sky130_fd_sc_hd__mux2_1
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27844_ _12298_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__clkbuf_1
X_20179_ registers\[48\]\[51\] registers\[49\]\[51\] registers\[50\]\[51\] registers\[51\]\[51\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__mux4_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24987_ _09646_ registers\[53\]\[63\] _10657_ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__mux2_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27775_ registers\[33\]\[36\] _10380_ _12255_ VGND VGND VPWR VPWR _12262_ sky130_fd_sc_hd__mux2_1
XFILLER_79_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29514_ _13207_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__clkbuf_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23938_ _10141_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26726_ _11678_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_700 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_898 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_711 _07303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_722 _07344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26657_ _10835_ registers\[41\]\[50\] _11641_ VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__mux2_1
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29445_ _13171_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_733 _07352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23869_ _10105_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_744 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_89_CLK sky130_fd_sc_hd__clkbuf_16
X_16410_ _14601_ _14913_ _14914_ _14611_ VGND VGND VPWR VPWR _14915_ sky130_fd_sc_hd__a22o_1
XANTENNA_755 _07385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25608_ registers\[48\]\[2\] _10309_ _11086_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__mux2_1
XANTENNA_766 _07639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17390_ _15830_ _15865_ _15866_ _15833_ VGND VGND VPWR VPWR _15867_ sky130_fd_sc_hd__a22o_1
X_29376_ _09819_ registers\[22\]\[60\] _13068_ VGND VGND VPWR VPWR _13135_ sky130_fd_sc_hd__mux2_1
XANTENNA_777 _08219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26588_ _11605_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_788 _08872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_799 _08936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16341_ _14847_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
X_28327_ _12552_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__clkbuf_1
X_25539_ registers\[4\]\[35\] _10378_ _11045_ VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__mux2_1
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19060_ _05496_ _05802_ _05803_ _05499_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__a22o_1
X_16272_ registers\[40\]\[6\] registers\[41\]\[6\] registers\[42\]\[6\] registers\[43\]\[6\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14780_ sky130_fd_sc_hd__mux4_1
X_28258_ registers\[2\]\[9\] _10323_ _12506_ VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__mux2_1
XFILLER_186_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18011_ _04779_ _04782_ _04611_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__o21ba_1
XFILLER_199_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27209_ _11963_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28189_ _11813_ registers\[30\]\[40\] _12479_ VGND VGND VPWR VPWR _12480_ sky130_fd_sc_hd__mux2_1
XFILLER_154_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30220_ _13579_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30151_ registers\[16\]\[43\] _13025_ _13539_ VGND VGND VPWR VPWR _13543_ sky130_fd_sc_hd__mux2_1
X_19962_ registers\[60\]\[45\] registers\[61\]\[45\] registers\[62\]\[45\] registers\[63\]\[45\]
+ _06648_ _06442_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__mux4_1
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_13_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18913_ registers\[4\]\[15\] registers\[5\]\[15\] registers\[6\]\[15\] registers\[7\]\[15\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__mux4_1
XTAP_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30082_ registers\[16\]\[10\] _12955_ _13506_ VGND VGND VPWR VPWR _13507_ sky130_fd_sc_hd__mux2_1
XTAP_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19893_ registers\[56\]\[43\] registers\[57\]\[43\] registers\[58\]\[43\] registers\[59\]\[43\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__mux4_1
XANTENNA_1110 _14564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1121 _14573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1132 _14607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33910_ clknet_leaf_336_CLK _02024_ VGND VGND VPWR VPWR registers\[38\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18844_ _05067_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__buf_4
XANTENNA_1143 _15041_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34890_ clknet_leaf_143_CLK _03004_ VGND VGND VPWR VPWR registers\[23\]\[60\] sky130_fd_sc_hd__dfxtp_1
XTAP_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1154 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1165 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1176 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1187 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33841_ clknet_leaf_381_CLK _01955_ VGND VGND VPWR VPWR registers\[3\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1198 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18775_ _05345_ _05525_ _05526_ _05348_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a22o_1
XFILLER_62_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15987_ _14500_ VGND VGND VPWR VPWR _14501_ sky130_fd_sc_hd__clkbuf_4
XTAP_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17726_ _14571_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__buf_4
X_33772_ clknet_leaf_325_CLK _01886_ VGND VGND VPWR VPWR registers\[40\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_30984_ _13981_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35511_ clknet_leaf_320_CLK _03625_ VGND VGND VPWR VPWR registers\[13\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32723_ clknet_leaf_72_CLK _00837_ VGND VGND VPWR VPWR registers\[56\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17657_ _04340_ _04437_ _04438_ _04343_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__a22o_1
X_16608_ _14504_ VGND VGND VPWR VPWR _15107_ sky130_fd_sc_hd__buf_4
X_35442_ clknet_leaf_380_CLK _03556_ VGND VGND VPWR VPWR registers\[14\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_23__f_CLK clknet_5_11_0_CLK VGND VGND VPWR VPWR clknet_6_23__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_32654_ clknet_leaf_74_CLK _00768_ VGND VGND VPWR VPWR registers\[57\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17588_ _04333_ _04370_ _04371_ _04338_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a22o_1
XFILLER_56_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31605_ registers\[63\]\[28\] net21 _14299_ VGND VGND VPWR VPWR _14308_ sky130_fd_sc_hd__mux2_1
X_19327_ _05747_ _06061_ _06062_ _05753_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__a22o_1
X_16539_ _14863_ _15038_ _15039_ _14867_ VGND VGND VPWR VPWR _15040_ sky130_fd_sc_hd__a22o_1
X_35373_ clknet_leaf_392_CLK _03487_ VGND VGND VPWR VPWR registers\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_32585_ clknet_leaf_161_CLK _00699_ VGND VGND VPWR VPWR registers\[5\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34324_ clknet_leaf_98_CLK _02438_ VGND VGND VPWR VPWR registers\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31536_ _14271_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19258_ _05755_ _05994_ _05995_ _05759_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__a22o_1
XFILLER_143_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18209_ registers\[28\]\[61\] registers\[29\]\[61\] registers\[30\]\[61\] registers\[31\]\[61\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__mux4_1
X_34255_ clknet_leaf_146_CLK _02369_ VGND VGND VPWR VPWR registers\[32\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31467_ _14235_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19189_ _05747_ _05927_ _05928_ _05753_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__a22o_1
XFILLER_191_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21220_ registers\[20\]\[15\] registers\[21\]\[15\] registers\[22\]\[15\] registers\[23\]\[15\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__mux4_1
X_33206_ clknet_leaf_319_CLK _01320_ VGND VGND VPWR VPWR registers\[4\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_30418_ _09778_ registers\[14\]\[41\] _13682_ VGND VGND VPWR VPWR _13684_ sky130_fd_sc_hd__mux2_1
X_34186_ clknet_leaf_156_CLK _02300_ VGND VGND VPWR VPWR registers\[34\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_31398_ registers\[7\]\[58\] net54 _14190_ VGND VGND VPWR VPWR _14199_ sky130_fd_sc_hd__mux2_1
XFILLER_145_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33137_ clknet_leaf_366_CLK _01251_ VGND VGND VPWR VPWR registers\[50\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_21151_ registers\[16\]\[13\] registers\[17\]\[13\] registers\[18\]\[13\] registers\[19\]\[13\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__mux4_1
XFILLER_172_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30349_ _13647_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20102_ _06812_ _06815_ _06504_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__o21ba_1
XFILLER_137_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21082_ _07732_ _07768_ _07769_ _07735_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__a22o_1
XFILLER_67_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33068_ clknet_leaf_379_CLK _01182_ VGND VGND VPWR VPWR registers\[51\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_20033_ _06433_ _06747_ _06748_ _06439_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__a22o_1
XFILLER_59_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24910_ _09569_ registers\[53\]\[26\] _10680_ VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32019_ clknet_leaf_182_CLK _00197_ VGND VGND VPWR VPWR registers\[62\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25890_ _10745_ registers\[46\]\[7\] _11230_ VGND VGND VPWR VPWR _11238_ sky130_fd_sc_hd__mux2_1
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24841_ _10650_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27560_ _12147_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24772_ _10614_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21984_ _08642_ _08645_ _08405_ _08406_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__o211a_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26511_ _11564_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35709_ clknet_leaf_300_CLK _03823_ VGND VGND VPWR VPWR registers\[10\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_23723_ _10016_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__buf_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _07373_ _07625_ _07626_ _07383_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__a22o_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27491_ _11792_ registers\[35\]\[30\] _12111_ VGND VGND VPWR VPWR _12112_ sky130_fd_sc_hd__mux2_1
XFILLER_163_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29230_ _13055_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26442_ _11528_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__clkbuf_1
X_23654_ _09990_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ registers\[28\]\[5\] registers\[29\]\[5\] registers\[30\]\[5\] registers\[31\]\[5\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__mux4_1
XFILLER_39_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22605_ registers\[40\]\[55\] registers\[41\]\[55\] registers\[42\]\[55\] registers\[43\]\[55\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__mux4_1
XFILLER_228_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29161_ registers\[23\]\[35\] _13008_ _12998_ VGND VGND VPWR VPWR _13009_ sky130_fd_sc_hd__mux2_1
X_26373_ _10823_ registers\[43\]\[44\] _11487_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23585_ _09942_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__buf_6
X_20797_ registers\[24\]\[3\] registers\[25\]\[3\] registers\[26\]\[3\] registers\[27\]\[3\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__mux4_1
X_28112_ _12439_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__clkbuf_1
X_25324_ _09867_ _10584_ VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__nor2_8
X_22536_ _09177_ _09182_ _09116_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__o21ba_1
XFILLER_128_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29092_ net5 VGND VGND VPWR VPWR _12962_ sky130_fd_sc_hd__buf_4
XFILLER_155_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28043_ _11803_ registers\[31\]\[35\] _12397_ VGND VGND VPWR VPWR _12403_ sky130_fd_sc_hd__mux2_1
X_25255_ _10899_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__clkbuf_1
X_22467_ _07398_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__clkbuf_2
XFILLER_183_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24206_ _10283_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21418_ _08092_ _08095_ _08054_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__o21ba_1
X_25186_ net60 VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__buf_2
X_22398_ _08805_ _09044_ _09047_ _08810_ VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__a22o_1
XFILLER_108_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24137_ _10247_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
X_21349_ _07991_ _08027_ _08028_ _07995_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__a22o_1
XFILLER_194_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29994_ _13460_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24068_ _10210_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
X_28945_ _12877_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23019_ net40 VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__clkbuf_4
XFILLER_235_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28876_ _11826_ registers\[25\]\[46\] _12834_ VGND VGND VPWR VPWR _12841_ sky130_fd_sc_hd__mux2_1
X_16890_ registers\[60\]\[23\] registers\[61\]\[23\] registers\[62\]\[23\] registers\[63\]\[23\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15381_ sky130_fd_sc_hd__mux4_1
X_27827_ registers\[33\]\[61\] _10432_ _12221_ VGND VGND VPWR VPWR _12289_ sky130_fd_sc_hd__mux2_1
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18560_ registers\[4\]\[5\] registers\[5\]\[5\] registers\[6\]\[5\] registers\[7\]\[5\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__mux4_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_24_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_24_0_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27758_ registers\[33\]\[28\] _10363_ _12244_ VGND VGND VPWR VPWR _12253_ sky130_fd_sc_hd__mux2_1
XFILLER_206_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17511_ registers\[20\]\[40\] registers\[21\]\[40\] registers\[22\]\[40\] registers\[23\]\[40\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__mux4_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26709_ registers\[40\]\[10\] _10325_ _11669_ VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__mux2_1
XFILLER_73_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18491_ _05120_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__buf_6
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27689_ _12216_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__clkbuf_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_530 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_884 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _14518_ VGND VGND VPWR VPWR _15917_ sky130_fd_sc_hd__buf_4
X_29428_ _09699_ registers\[21\]\[20\] _13162_ VGND VGND VPWR VPWR _13163_ sky130_fd_sc_hd__mux2_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_552 _04675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_563 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_2_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_574 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_585 _05067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_596 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29359_ _13126_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__clkbuf_1
X_17373_ _14571_ VGND VGND VPWR VPWR _15850_ sky130_fd_sc_hd__buf_4
XFILLER_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19112_ registers\[40\]\[21\] registers\[41\]\[21\] registers\[42\]\[21\] registers\[43\]\[21\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__mux4_1
X_16324_ _14540_ _14829_ _14830_ _14551_ VGND VGND VPWR VPWR _14831_ sky130_fd_sc_hd__a22o_1
XFILLER_13_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32370_ clknet_leaf_356_CLK _00484_ VGND VGND VPWR VPWR registers\[61\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16255_ _14504_ VGND VGND VPWR VPWR _14764_ sky130_fd_sc_hd__buf_4
X_31321_ registers\[7\]\[21\] net14 _14157_ VGND VGND VPWR VPWR _14159_ sky130_fd_sc_hd__mux2_1
X_19043_ _05783_ _05786_ _05475_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__o21ba_1
XFILLER_127_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31252_ _14122_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34040_ clknet_leaf_337_CLK _02154_ VGND VGND VPWR VPWR registers\[36\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_16186_ _14540_ _14695_ _14696_ _14551_ VGND VGND VPWR VPWR _14697_ sky130_fd_sc_hd__a22o_1
Xoutput206 net206 VGND VGND VPWR VPWR D2[57] sky130_fd_sc_hd__buf_2
XFILLER_127_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 net217 VGND VGND VPWR VPWR D2[9] sky130_fd_sc_hd__buf_2
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30203_ _13570_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput228 net228 VGND VGND VPWR VPWR D3[19] sky130_fd_sc_hd__buf_2
X_31183_ _14063_ VGND VGND VPWR VPWR _14086_ sky130_fd_sc_hd__buf_4
XFILLER_142_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput239 net239 VGND VGND VPWR VPWR D3[29] sky130_fd_sc_hd__buf_2
XFILLER_5_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30134_ registers\[16\]\[35\] _13008_ _13528_ VGND VGND VPWR VPWR _13534_ sky130_fd_sc_hd__mux2_1
XFILLER_138_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19945_ _06525_ _06662_ _06663_ _06528_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__a22o_1
XFILLER_218_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35991_ clknet_leaf_61_CLK _04105_ VGND VGND VPWR VPWR registers\[63\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30065_ registers\[16\]\[2\] _12939_ _13495_ VGND VGND VPWR VPWR _13498_ sky130_fd_sc_hd__mux2_1
X_34942_ clknet_leaf_187_CLK _03056_ VGND VGND VPWR VPWR registers\[22\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_19876_ registers\[16\]\[42\] registers\[17\]\[42\] registers\[18\]\[42\] registers\[19\]\[42\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__mux4_1
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18827_ registers\[40\]\[13\] registers\[41\]\[13\] registers\[42\]\[13\] registers\[43\]\[13\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__mux4_1
X_34873_ clknet_leaf_309_CLK _02987_ VGND VGND VPWR VPWR registers\[23\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33824_ clknet_leaf_486_CLK _01938_ VGND VGND VPWR VPWR registers\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_18758_ _05510_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17709_ _04486_ _04487_ _04488_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a22o_1
XFILLER_208_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33755_ clknet_leaf_25_CLK _01869_ VGND VGND VPWR VPWR registers\[40\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_18689_ _05204_ _05441_ _05442_ _05207_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__a22o_1
X_30967_ _13972_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20720_ registers\[8\]\[1\] registers\[9\]\[1\] registers\[10\]\[1\] registers\[11\]\[1\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__mux4_1
X_32706_ clknet_leaf_263_CLK _00820_ VGND VGND VPWR VPWR registers\[57\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_33686_ clknet_leaf_126_CLK _01800_ VGND VGND VPWR VPWR registers\[41\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30898_ _13936_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35425_ clknet_leaf_482_CLK _03539_ VGND VGND VPWR VPWR registers\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20651_ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__clkbuf_4
X_32637_ clknet_leaf_289_CLK _00751_ VGND VGND VPWR VPWR registers\[58\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35356_ clknet_leaf_477_CLK _03470_ VGND VGND VPWR VPWR registers\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_23370_ _09838_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
X_20582_ _07280_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__buf_12
XFILLER_149_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32568_ clknet_leaf_314_CLK _00682_ VGND VGND VPWR VPWR registers\[5\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34307_ clknet_leaf_250_CLK _02421_ VGND VGND VPWR VPWR registers\[32\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_22321_ _08973_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_2
XFILLER_109_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31519_ _09800_ registers\[6\]\[51\] _14261_ VGND VGND VPWR VPWR _14263_ sky130_fd_sc_hd__mux2_1
XFILLER_191_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35287_ clknet_leaf_91_CLK _03401_ VGND VGND VPWR VPWR registers\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32499_ clknet_leaf_357_CLK _00613_ VGND VGND VPWR VPWR registers\[60\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_25040_ _10763_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
X_34238_ clknet_leaf_268_CLK _02352_ VGND VGND VPWR VPWR registers\[33\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_22252_ registers\[40\]\[45\] registers\[41\]\[45\] registers\[42\]\[45\] registers\[43\]\[45\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__mux4_1
XFILLER_129_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21203_ registers\[60\]\[15\] registers\[61\]\[15\] registers\[62\]\[15\] registers\[63\]\[15\]
+ _07855_ _07649_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__mux4_1
XFILLER_145_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22183_ _08834_ _08839_ _08773_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__o21ba_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34169_ clknet_leaf_336_CLK _02283_ VGND VGND VPWR VPWR registers\[34\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21134_ registers\[56\]\[13\] registers\[57\]\[13\] registers\[58\]\[13\] registers\[59\]\[13\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__mux4_1
XFILLER_156_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26991_ _11843_ registers\[3\]\[54\] _11835_ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__mux2_1
XFILLER_120_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28730_ _12764_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21065_ _07749_ _07752_ _07711_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__o21ba_1
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25942_ _11265_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20016_ registers\[28\]\[46\] registers\[29\]\[46\] registers\[30\]\[46\] registers\[31\]\[46\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__mux4_1
XFILLER_48_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25873_ _11228_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
X_28661_ _11746_ registers\[26\]\[8\] _12719_ VGND VGND VPWR VPWR _12728_ sky130_fd_sc_hd__mux2_1
XFILLER_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24824_ _10641_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27612_ _12176_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28592_ _12691_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27543_ _11845_ registers\[35\]\[55\] _12133_ VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__mux2_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24755_ _10605_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
X_21967_ _08600_ _08609_ _08620_ _08629_ VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__or4_1
XFILLER_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23706_ _10019_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _07604_ _07609_ _07310_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__o21ba_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27474_ _11776_ registers\[35\]\[22\] _12100_ VGND VGND VPWR VPWR _12103_ sky130_fd_sc_hd__mux2_1
X_24686_ _09617_ registers\[55\]\[49\] _10558_ VGND VGND VPWR VPWR _10568_ sky130_fd_sc_hd__mux2_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21898_ _08562_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__buf_6
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29213_ net48 VGND VGND VPWR VPWR _13044_ sky130_fd_sc_hd__clkbuf_4
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26425_ _11519_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23637_ _09981_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20849_ _07313_ _07541_ _07542_ _07322_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__a22o_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29144_ net24 VGND VGND VPWR VPWR _12997_ sky130_fd_sc_hd__buf_2
X_26356_ _10806_ registers\[43\]\[36\] _11476_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23568_ _09945_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25307_ _10926_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22519_ _09020_ _09164_ _09165_ _09024_ VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__a22o_1
X_26287_ _10737_ registers\[43\]\[3\] _11443_ VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__mux2_1
X_29075_ _12950_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__clkbuf_1
X_23499_ _09586_ registers\[19\]\[34\] _09903_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__mux2_1
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _14553_ VGND VGND VPWR VPWR _14554_ sky130_fd_sc_hd__buf_2
XFILLER_183_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28026_ _11786_ registers\[31\]\[27\] _12386_ VGND VGND VPWR VPWR _12394_ sky130_fd_sc_hd__mux2_1
X_25238_ _10890_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25169_ _10850_ registers\[52\]\[57\] _10836_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__mux2_1
X_17991_ registers\[4\]\[54\] registers\[5\]\[54\] registers\[6\]\[54\] registers\[7\]\[54\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__mux4_1
X_29977_ _13451_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19730_ _06379_ _06451_ _06454_ _06382_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__a22o_1
X_28928_ _12868_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__clkbuf_1
X_16942_ _15295_ _15430_ _15431_ _15300_ VGND VGND VPWR VPWR _15432_ sky130_fd_sc_hd__a22o_1
XFILLER_237_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19661_ registers\[16\]\[36\] registers\[17\]\[36\] registers\[18\]\[36\] registers\[19\]\[36\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__mux4_1
XFILLER_81_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16873_ _14603_ VGND VGND VPWR VPWR _15365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28859_ _11809_ registers\[25\]\[38\] _12823_ VGND VGND VPWR VPWR _12832_ sky130_fd_sc_hd__mux2_1
X_18612_ _05197_ _05366_ _05367_ _05202_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__a22o_1
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _06182_ _06319_ _06320_ _06185_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__a22o_1
X_31870_ _14447_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__clkbuf_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ registers\[44\]\[5\] registers\[45\]\[5\] registers\[46\]\[5\] registers\[47\]\[5\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__mux4_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30821_ _09775_ registers\[11\]\[40\] _13895_ VGND VGND VPWR VPWR _13896_ sky130_fd_sc_hd__mux2_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33540_ clknet_leaf_251_CLK _01654_ VGND VGND VPWR VPWR registers\[44\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18474_ registers\[40\]\[3\] registers\[41\]\[3\] registers\[42\]\[3\] registers\[43\]\[3\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__mux4_1
X_30752_ _13859_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_360 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_382 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ _15825_ _15899_ _15900_ _15828_ VGND VGND VPWR VPWR _15901_ sky130_fd_sc_hd__a22o_1
XANTENNA_393 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33471_ clknet_leaf_273_CLK _01585_ VGND VGND VPWR VPWR registers\[45\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30683_ registers\[12\]\[39\] _13016_ _13813_ VGND VGND VPWR VPWR _13823_ sky130_fd_sc_hd__mux2_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35210_ clknet_leaf_149_CLK _03324_ VGND VGND VPWR VPWR registers\[18\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32422_ clknet_leaf_455_CLK _00536_ VGND VGND VPWR VPWR registers\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_36190_ clknet_leaf_91_CLK _00071_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_1
X_17356_ _15830_ _15831_ _15832_ _15833_ VGND VGND VPWR VPWR _15834_ sky130_fd_sc_hd__a22o_1
XFILLER_119_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35141_ clknet_leaf_228_CLK _03255_ VGND VGND VPWR VPWR registers\[1\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_16307_ _14811_ _14814_ _14614_ VGND VGND VPWR VPWR _14815_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32353_ clknet_leaf_44_CLK _00467_ VGND VGND VPWR VPWR registers\[61\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_17287_ _15763_ _15766_ _15631_ VGND VGND VPWR VPWR _15767_ sky130_fd_sc_hd__o21ba_1
XFILLER_179_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19026_ registers\[24\]\[18\] registers\[25\]\[18\] registers\[26\]\[18\] registers\[27\]\[18\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__mux4_1
X_31304_ registers\[7\]\[13\] net5 _14146_ VGND VGND VPWR VPWR _14150_ sky130_fd_sc_hd__mux2_1
X_35072_ clknet_leaf_203_CLK _03186_ VGND VGND VPWR VPWR registers\[20\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_16238_ _14722_ _14731_ _14738_ _14747_ VGND VGND VPWR VPWR _14748_ sky130_fd_sc_hd__or4_1
X_32284_ clknet_leaf_5_CLK _00398_ VGND VGND VPWR VPWR registers\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34023_ clknet_leaf_434_CLK _02137_ VGND VGND VPWR VPWR registers\[36\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_31235_ _14113_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__clkbuf_1
X_16169_ registers\[20\]\[2\] registers\[21\]\[2\] registers\[22\]\[2\] registers\[23\]\[2\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14681_ sky130_fd_sc_hd__mux4_1
XFILLER_173_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31166_ _14077_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19928_ _06433_ _06645_ _06646_ _06439_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__a22o_1
X_30117_ registers\[16\]\[27\] _12991_ _13517_ VGND VGND VPWR VPWR _13525_ sky130_fd_sc_hd__mux2_1
X_35974_ clknet_leaf_210_CLK _04088_ VGND VGND VPWR VPWR registers\[6\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_31097_ registers\[0\]\[43\] _13025_ _14037_ VGND VGND VPWR VPWR _14041_ sky130_fd_sc_hd__mux2_1
XFILLER_60_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30048_ _13488_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__clkbuf_1
X_34925_ clknet_leaf_402_CLK _03039_ VGND VGND VPWR VPWR registers\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_19859_ _06576_ _06577_ _06578_ _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__a22o_1
XFILLER_112_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22870_ registers\[20\]\[63\] registers\[21\]\[63\] registers\[22\]\[63\] registers\[23\]\[63\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__mux4_1
XFILLER_151_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34856_ clknet_leaf_454_CLK _02970_ VGND VGND VPWR VPWR registers\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33807_ clknet_leaf_135_CLK _01921_ VGND VGND VPWR VPWR registers\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_21821_ _08484_ _08487_ _08416_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__o21ba_1
XFILLER_71_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34787_ clknet_leaf_446_CLK _02901_ VGND VGND VPWR VPWR registers\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_31999_ clknet_leaf_29_CLK _00171_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_1
XFILLER_70_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24540_ _09609_ registers\[56\]\[45\] _10484_ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__mux2_1
X_33738_ clknet_leaf_161_CLK _01852_ VGND VGND VPWR VPWR registers\[41\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_21752_ _07382_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20703_ _07401_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
X_24471_ _09540_ registers\[56\]\[12\] _10451_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__mux2_1
XFILLER_52_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33669_ clknet_leaf_250_CLK _01783_ VGND VGND VPWR VPWR registers\[42\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_21683_ registers\[20\]\[28\] registers\[21\]\[28\] registers\[22\]\[28\] registers\[23\]\[28\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__mux4_1
X_26210_ _11406_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
X_35408_ clknet_leaf_138_CLK _03522_ VGND VGND VPWR VPWR registers\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_23422_ _09865_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__clkbuf_1
X_20634_ _07280_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__buf_12
XFILLER_71_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27190_ _11953_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26141_ _11369_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
X_35339_ clknet_leaf_149_CLK _03453_ VGND VGND VPWR VPWR registers\[16\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23353_ registers\[39\]\[30\] _09753_ _09829_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__mux2_1
X_20565_ _07261_ _07264_ _05133_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__o21ba_1
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22304_ _08953_ _08954_ _08955_ _08956_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__a22o_1
X_26072_ _11333_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23284_ registers\[9\]\[44\] _09784_ _09776_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__mux2_1
X_20496_ registers\[52\]\[61\] registers\[53\]\[61\] registers\[54\]\[61\] registers\[55\]\[61\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__mux4_1
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29900_ registers\[18\]\[52\] _13044_ _13408_ VGND VGND VPWR VPWR _13411_ sky130_fd_sc_hd__mux2_1
XFILLER_146_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25023_ _10730_ VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__buf_4
XFILLER_192_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22235_ registers\[0\]\[44\] registers\[1\]\[44\] registers\[2\]\[44\] registers\[3\]\[44\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__mux4_1
XFILLER_161_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29831_ _13374_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__clkbuf_1
X_22166_ _08677_ _08821_ _08822_ _08681_ VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__a22o_1
XTAP_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1709 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21117_ registers\[16\]\[12\] registers\[17\]\[12\] registers\[18\]\[12\] registers\[19\]\[12\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__mux4_1
X_29762_ _13338_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_1452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26974_ net44 VGND VGND VPWR VPWR _11832_ sky130_fd_sc_hd__clkbuf_4
X_22097_ registers\[12\]\[40\] registers\[13\]\[40\] registers\[14\]\[40\] registers\[15\]\[40\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__mux4_1
XTAP_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28713_ _12755_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__clkbuf_1
X_25925_ _11256_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
X_21048_ _07385_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__buf_4
X_29693_ registers\[1\]\[18\] _12972_ _13293_ VGND VGND VPWR VPWR _13302_ sky130_fd_sc_hd__mux2_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28644_ _12718_ VGND VGND VPWR VPWR _12719_ sky130_fd_sc_hd__buf_4
XFILLER_86_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25856_ _10846_ registers\[47\]\[55\] _11214_ VGND VGND VPWR VPWR _11220_ sky130_fd_sc_hd__mux2_1
XFILLER_74_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24807_ _09601_ registers\[54\]\[41\] _10631_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__mux2_1
X_28575_ _11795_ registers\[27\]\[31\] _12681_ VGND VGND VPWR VPWR _12683_ sky130_fd_sc_hd__mux2_1
X_25787_ _10777_ registers\[47\]\[22\] _11181_ VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__mux2_1
XFILLER_43_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22999_ _09595_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_27526_ _11828_ registers\[35\]\[47\] _12122_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__mux2_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24738_ _10596_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27457_ _11759_ registers\[35\]\[14\] _12089_ VGND VGND VPWR VPWR _12094_ sky130_fd_sc_hd__mux2_1
X_24669_ _10559_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17210_ _15541_ _15690_ _15691_ _15547_ VGND VGND VPWR VPWR _15692_ sky130_fd_sc_hd__a22o_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26408_ _10858_ registers\[43\]\[61\] _11442_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18190_ _04683_ _04954_ _04955_ _04686_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__a22o_1
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27388_ _12057_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17141_ _14564_ VGND VGND VPWR VPWR _15625_ sky130_fd_sc_hd__clkbuf_4
X_29127_ registers\[23\]\[24\] _12985_ _12977_ VGND VGND VPWR VPWR _12986_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26339_ _10789_ registers\[43\]\[28\] _11465_ VGND VGND VPWR VPWR _11474_ sky130_fd_sc_hd__mux2_1
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17072_ _15482_ _15556_ _15557_ _15485_ VGND VGND VPWR VPWR _15558_ sky130_fd_sc_hd__a22o_1
X_29058_ net23 VGND VGND VPWR VPWR _12939_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16023_ _14500_ VGND VGND VPWR VPWR _14537_ sky130_fd_sc_hd__buf_2
X_28009_ _11769_ registers\[31\]\[19\] _12375_ VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__mux2_1
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31020_ _14000_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17974_ registers\[44\]\[54\] registers\[45\]\[54\] registers\[46\]\[54\] registers\[47\]\[54\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__mux4_1
X_19713_ registers\[48\]\[38\] registers\[49\]\[38\] registers\[50\]\[38\] registers\[51\]\[38\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__mux4_1
XFILLER_111_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16925_ registers\[52\]\[24\] registers\[53\]\[24\] registers\[54\]\[24\] registers\[55\]\[24\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15415_ sky130_fd_sc_hd__mux4_1
XFILLER_66_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32971_ clknet_leaf_166_CLK _01085_ VGND VGND VPWR VPWR registers\[53\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_293_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_293_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34710_ clknet_leaf_88_CLK _02824_ VGND VGND VPWR VPWR registers\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31922_ _09797_ registers\[49\]\[50\] _14474_ VGND VGND VPWR VPWR _14475_ sky130_fd_sc_hd__mux2_1
X_19644_ registers\[52\]\[36\] registers\[53\]\[36\] registers\[54\]\[36\] registers\[55\]\[36\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__mux4_1
X_35690_ clknet_leaf_399_CLK _03804_ VGND VGND VPWR VPWR registers\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_16856_ registers\[48\]\[22\] registers\[49\]\[22\] registers\[50\]\[22\] registers\[51\]\[22\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15348_ sky130_fd_sc_hd__mux4_1
XFILLER_238_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34641_ clknet_leaf_117_CLK _02755_ VGND VGND VPWR VPWR registers\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_19575_ _06090_ _06302_ _06303_ _06096_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__a22o_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31853_ _14438_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__clkbuf_1
X_16787_ _14562_ VGND VGND VPWR VPWR _15281_ sky130_fd_sc_hd__buf_6
XFILLER_4_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18526_ registers\[4\]\[4\] registers\[5\]\[4\] registers\[6\]\[4\] registers\[7\]\[4\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__mux4_1
X_30804_ _09758_ registers\[11\]\[32\] _13884_ VGND VGND VPWR VPWR _13887_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34572_ clknet_leaf_141_CLK _02686_ VGND VGND VPWR VPWR registers\[28\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31784_ registers\[59\]\[49\] net44 _14392_ VGND VGND VPWR VPWR _14402_ sky130_fd_sc_hd__mux2_1
XFILLER_221_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33523_ clknet_leaf_346_CLK _01637_ VGND VGND VPWR VPWR registers\[44\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_30735_ _13636_ _09868_ VGND VGND VPWR VPWR _13850_ sky130_fd_sc_hd__nand2_8
X_18457_ registers\[0\]\[2\] registers\[1\]\[2\] registers\[2\]\[2\] registers\[3\]\[2\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__mux4_1
XFILLER_205_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_190 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_222_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17408_ _14527_ VGND VGND VPWR VPWR _15884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_222_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33454_ clknet_leaf_360_CLK _01568_ VGND VGND VPWR VPWR registers\[45\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_18388_ _05141_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__buf_6
X_30666_ _13814_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32405_ clknet_leaf_95_CLK _00519_ VGND VGND VPWR VPWR registers\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_36173_ clknet_leaf_170_CLK _04287_ VGND VGND VPWR VPWR registers\[49\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_17339_ registers\[48\]\[36\] registers\[49\]\[36\] registers\[50\]\[36\] registers\[51\]\[36\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15817_ sky130_fd_sc_hd__mux4_1
X_33385_ clknet_leaf_60_CLK _01499_ VGND VGND VPWR VPWR registers\[46\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_30597_ _13777_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35124_ clknet_leaf_414_CLK _03238_ VGND VGND VPWR VPWR registers\[1\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_20350_ registers\[0\]\[56\] registers\[1\]\[56\] registers\[2\]\[56\] registers\[3\]\[56\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__mux4_1
X_32336_ clknet_leaf_175_CLK _00450_ VGND VGND VPWR VPWR registers\[61\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19009_ _05747_ _05749_ _05752_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__a22o_1
X_35055_ clknet_leaf_395_CLK _03169_ VGND VGND VPWR VPWR registers\[20\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_32267_ clknet_leaf_165_CLK _00381_ VGND VGND VPWR VPWR registers\[39\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_20281_ _06776_ _06988_ _06989_ _06782_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__a22o_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34006_ clknet_leaf_120_CLK _02120_ VGND VGND VPWR VPWR registers\[36\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_22020_ _07301_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__clkbuf_4
X_31218_ _14104_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32198_ clknet_leaf_391_CLK _00312_ VGND VGND VPWR VPWR registers\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31149_ _14068_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__clkbuf_1
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23971_ _10158_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35957_ clknet_leaf_322_CLK _04071_ VGND VGND VPWR VPWR registers\[6\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_284_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_284_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25710_ _11142_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
X_22922_ _09543_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26690_ registers\[40\]\[1\] _10307_ _11658_ VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__mux2_1
X_34908_ clknet_leaf_492_CLK _03022_ VGND VGND VPWR VPWR registers\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_35888_ clknet_leaf_374_CLK _04002_ VGND VGND VPWR VPWR registers\[7\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22853_ registers\[48\]\[63\] registers\[49\]\[63\] registers\[50\]\[63\] registers\[51\]\[63\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__mux4_1
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25641_ registers\[48\]\[18\] _10342_ _11097_ VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34839_ clknet_leaf_99_CLK _02953_ VGND VGND VPWR VPWR registers\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21804_ registers\[36\]\[32\] registers\[37\]\[32\] registers\[38\]\[32\] registers\[39\]\[32\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__mux4_1
X_28360_ _12569_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__clkbuf_1
X_25572_ _11068_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
X_22784_ _09422_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27311_ registers\[36\]\[9\] _10323_ _12007_ VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__mux2_1
XFILLER_212_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24523_ _09592_ registers\[56\]\[37\] _10473_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__mux2_1
X_21735_ _08334_ _08402_ _08403_ _08338_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__a22o_1
XFILLER_213_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28291_ _12533_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_835 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24454_ _09523_ registers\[56\]\[4\] _10440_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__mux2_1
X_27242_ _11813_ registers\[37\]\[40\] _11980_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__mux2_1
X_21666_ registers\[52\]\[28\] registers\[53\]\[28\] registers\[54\]\[28\] registers\[55\]\[28\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__mux4_1
XFILLER_71_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23405_ registers\[39\]\[55\] _09808_ _09851_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27173_ _11944_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_1
X_20617_ _07280_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__buf_12
X_24385_ net40 VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__clkbuf_4
XFILLER_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21597_ _07352_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__buf_4
X_26124_ _10844_ registers\[45\]\[54\] _11356_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__mux2_1
X_23336_ net57 VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__clkbuf_4
X_20548_ registers\[44\]\[63\] registers\[45\]\[63\] registers\[46\]\[63\] registers\[47\]\[63\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__mux4_1
XFILLER_193_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26055_ _10775_ registers\[45\]\[21\] _11323_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__mux2_1
X_23267_ net33 VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__clkbuf_4
X_20479_ registers\[28\]\[60\] registers\[29\]\[60\] registers\[30\]\[60\] registers\[31\]\[60\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__mux4_1
XFILLER_197_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25006_ _10740_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
X_22218_ registers\[40\]\[44\] registers\[41\]\[44\] registers\[42\]\[44\] registers\[43\]\[44\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__mux4_1
XFILLER_234_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23198_ _09729_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1506 _07382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1517 _08841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29814_ registers\[18\]\[11\] _12958_ _13364_ VGND VGND VPWR VPWR _13366_ sky130_fd_sc_hd__mux2_1
XTAP_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22149_ _07278_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__buf_4
XTAP_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1528 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1539 _09793_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29745_ _13329_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26957_ _11820_ registers\[3\]\[43\] _11814_ VGND VGND VPWR VPWR _11821_ sky130_fd_sc_hd__mux2_1
XTAP_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_275_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_275_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16710_ _14539_ VGND VGND VPWR VPWR _15206_ sky130_fd_sc_hd__clkbuf_4
XFILLER_248_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25908_ _11247_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17690_ _04467_ _04470_ _15955_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__o21ba_1
X_29676_ _13281_ VGND VGND VPWR VPWR _13293_ sky130_fd_sc_hd__buf_4
XFILLER_48_968 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26888_ net14 VGND VGND VPWR VPWR _11774_ sky130_fd_sc_hd__clkbuf_4
X_28627_ _11847_ registers\[27\]\[56\] _12703_ VGND VGND VPWR VPWR _12710_ sky130_fd_sc_hd__mux2_1
X_16641_ _14490_ VGND VGND VPWR VPWR _15139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25839_ _10829_ registers\[47\]\[47\] _11203_ VGND VGND VPWR VPWR _11211_ sky130_fd_sc_hd__mux2_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19360_ registers\[48\]\[28\] registers\[49\]\[28\] registers\[50\]\[28\] registers\[51\]\[28\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__mux4_1
X_16572_ registers\[52\]\[14\] registers\[53\]\[14\] registers\[54\]\[14\] registers\[55\]\[14\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _15072_ sky130_fd_sc_hd__mux4_1
X_28558_ _11778_ registers\[27\]\[23\] _12670_ VGND VGND VPWR VPWR _12674_ sky130_fd_sc_hd__mux2_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18311_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__buf_2
XFILLER_16_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27509_ _11811_ registers\[35\]\[39\] _12111_ VGND VGND VPWR VPWR _12121_ sky130_fd_sc_hd__mux2_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19291_ registers\[52\]\[26\] registers\[53\]\[26\] registers\[54\]\[26\] registers\[55\]\[26\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__mux4_1
X_28489_ _12637_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18242_ _05003_ _05006_ _14613_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__o21ba_1
XFILLER_203_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30520_ _13737_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__clkbuf_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30451_ _09813_ registers\[14\]\[57\] _13693_ VGND VGND VPWR VPWR _13701_ sky130_fd_sc_hd__mux2_1
X_18173_ registers\[4\]\[60\] registers\[5\]\[60\] registers\[6\]\[60\] registers\[7\]\[60\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__mux4_1
XFILLER_50_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17124_ _14548_ VGND VGND VPWR VPWR _15608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33170_ clknet_leaf_77_CLK _01284_ VGND VGND VPWR VPWR registers\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30382_ _09740_ registers\[14\]\[24\] _13660_ VGND VGND VPWR VPWR _13665_ sky130_fd_sc_hd__mux2_1
XFILLER_144_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32121_ clknet_leaf_393_CLK _00037_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17055_ _14527_ VGND VGND VPWR VPWR _15541_ sky130_fd_sc_hd__buf_4
X_16006_ _14495_ VGND VGND VPWR VPWR _14520_ sky130_fd_sc_hd__buf_12
XFILLER_125_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32052_ clknet_leaf_325_CLK _00230_ VGND VGND VPWR VPWR registers\[62\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31003_ registers\[10\]\[63\] _13066_ _13921_ VGND VGND VPWR VPWR _13991_ sky130_fd_sc_hd__mux2_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35811_ clknet_leaf_466_CLK _03925_ VGND VGND VPWR VPWR registers\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17957_ _14520_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__buf_4
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_266_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_266_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35742_ clknet_leaf_479_CLK _03856_ VGND VGND VPWR VPWR registers\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_16908_ _15295_ _15397_ _15398_ _15300_ VGND VGND VPWR VPWR _15399_ sky130_fd_sc_hd__a22o_1
XFILLER_238_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32954_ clknet_leaf_286_CLK _01068_ VGND VGND VPWR VPWR registers\[53\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_17888_ registers\[12\]\[51\] registers\[13\]\[51\] registers\[14\]\[51\] registers\[15\]\[51\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__mux4_1
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31905_ _09780_ registers\[49\]\[42\] _14463_ VGND VGND VPWR VPWR _14466_ sky130_fd_sc_hd__mux2_1
X_19627_ _06187_ _06353_ _06354_ _06192_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__a22o_1
X_16839_ _15328_ _15331_ _15302_ VGND VGND VPWR VPWR _15332_ sky130_fd_sc_hd__o21ba_1
X_35673_ clknet_leaf_12_CLK _03787_ VGND VGND VPWR VPWR registers\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32885_ clknet_leaf_352_CLK _00999_ VGND VGND VPWR VPWR registers\[54\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34624_ clknet_leaf_224_CLK _02738_ VGND VGND VPWR VPWR registers\[27\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31836_ _14429_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__clkbuf_1
X_19558_ _06182_ _06286_ _06287_ _06185_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__a22o_1
XFILLER_59_1262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18509_ registers\[44\]\[4\] registers\[45\]\[4\] registers\[46\]\[4\] registers\[47\]\[4\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__mux4_1
X_34555_ clknet_leaf_184_CLK _02669_ VGND VGND VPWR VPWR registers\[28\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_19489_ registers\[28\]\[31\] registers\[29\]\[31\] registers\[30\]\[31\] registers\[31\]\[31\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux4_1
X_31767_ _14393_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33506_ clknet_leaf_58_CLK _01620_ VGND VGND VPWR VPWR registers\[44\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_21520_ registers\[56\]\[24\] registers\[57\]\[24\] registers\[58\]\[24\] registers\[59\]\[24\]
+ _08194_ _07984_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__mux4_1
X_30718_ _13841_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__clkbuf_1
X_34486_ clknet_leaf_318_CLK _02600_ VGND VGND VPWR VPWR registers\[2\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_31698_ registers\[59\]\[8\] net63 _14348_ VGND VGND VPWR VPWR _14357_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36225_ clknet_leaf_117_CLK _00110_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33437_ clknet_leaf_30_CLK _01551_ VGND VGND VPWR VPWR registers\[45\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_21451_ registers\[36\]\[22\] registers\[37\]\[22\] registers\[38\]\[22\] registers\[39\]\[22\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__mux4_1
X_30649_ _13805_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__clkbuf_1
X_20402_ registers\[56\]\[58\] registers\[57\]\[58\] registers\[58\]\[58\] registers\[59\]\[58\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__mux4_1
XFILLER_175_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36156_ clknet_leaf_282_CLK _04270_ VGND VGND VPWR VPWR registers\[49\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_24170_ _10264_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
X_33368_ clknet_leaf_31_CLK _01482_ VGND VGND VPWR VPWR registers\[46\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_21382_ _07991_ _08059_ _08060_ _07995_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__a22o_1
XFILLER_190_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35107_ clknet_leaf_471_CLK _03221_ VGND VGND VPWR VPWR registers\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_23121_ net3 VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__buf_6
X_20333_ _07019_ _07026_ _07033_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__or4_2
X_32319_ clknet_leaf_196_CLK _00433_ VGND VGND VPWR VPWR registers\[19\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_36087_ clknet_leaf_328_CLK _04201_ VGND VGND VPWR VPWR registers\[59\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_33299_ clknet_leaf_125_CLK _01413_ VGND VGND VPWR VPWR registers\[47\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23052_ _09631_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_1
X_35038_ clknet_leaf_490_CLK _03152_ VGND VGND VPWR VPWR registers\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_20264_ _06868_ _06972_ _06973_ _06871_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a22o_1
XTAP_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22003_ _08462_ _08662_ _08663_ _08467_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__a22o_1
XTAP_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27860_ registers\[32\]\[12\] _10330_ _12304_ VGND VGND VPWR VPWR _12307_ sky130_fd_sc_hd__mux2_1
X_20195_ registers\[28\]\[51\] registers\[29\]\[51\] registers\[30\]\[51\] registers\[31\]\[51\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__mux4_1
XTAP_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26811_ registers\[40\]\[59\] _10428_ _11713_ VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__mux2_1
XTAP_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27791_ _12270_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_257_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_257_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29530_ _13216_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26742_ registers\[40\]\[26\] _10359_ _11680_ VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__mux2_1
XFILLER_229_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23954_ _09630_ registers\[60\]\[55\] _10144_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__mux2_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22905_ _09531_ registers\[62\]\[8\] _09515_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__mux2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29461_ _09766_ registers\[21\]\[36\] _13173_ VGND VGND VPWR VPWR _13180_ sky130_fd_sc_hd__mux2_1
X_26673_ _10852_ registers\[41\]\[58\] _11641_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__mux2_1
X_23885_ _09561_ registers\[60\]\[22\] _10111_ VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__mux2_1
XFILLER_244_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_904 _09662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_915 _09708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28412_ _11767_ registers\[28\]\[18\] _12588_ VGND VGND VPWR VPWR _12597_ sky130_fd_sc_hd__mux2_1
X_22836_ registers\[24\]\[62\] registers\[25\]\[62\] registers\[26\]\[62\] registers\[27\]\[62\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__mux4_1
XANTENNA_926 _09817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25624_ _11085_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__buf_4
X_29392_ _09664_ registers\[21\]\[3\] _13140_ VGND VGND VPWR VPWR _13144_ sky130_fd_sc_hd__mux2_1
XANTENNA_937 _10232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_948 _10405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_959 _10814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_213_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28343_ _12560_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22767_ _07385_ _09404_ _09405_ _07395_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__a22o_1
X_25555_ _11059_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__clkbuf_1
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21718_ _08366_ _08373_ _08380_ _08387_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__or4_4
X_24506_ _09575_ registers\[56\]\[29\] _10462_ VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__mux2_1
XFILLER_197_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28274_ _12524_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25486_ _11011_ VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__buf_4
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22698_ registers\[44\]\[58\] registers\[45\]\[58\] registers\[46\]\[58\] registers\[47\]\[58\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__mux4_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27225_ _11797_ registers\[37\]\[32\] _11969_ VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__mux2_1
X_24437_ net59 VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21649_ registers\[32\]\[28\] registers\[33\]\[28\] registers\[34\]\[28\] registers\[35\]\[28\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__mux4_1
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27156_ _11863_ _10015_ VGND VGND VPWR VPWR _11935_ sky130_fd_sc_hd__nand2_8
XFILLER_138_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24368_ _10387_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_90 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23319_ net51 VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__buf_4
X_26107_ _10827_ registers\[45\]\[46\] _11345_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__mux2_1
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27087_ _11899_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_1
X_24299_ registers\[57\]\[17\] _10340_ _10326_ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__mux2_1
XFILLER_192_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26038_ _10758_ registers\[45\]\[13\] _11312_ VGND VGND VPWR VPWR _11316_ sky130_fd_sc_hd__mux2_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1303 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18860_ registers\[32\]\[14\] registers\[33\]\[14\] registers\[34\]\[14\] registers\[35\]\[14\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__mux4_1
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1314 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1325 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1336 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17811_ registers\[0\]\[49\] registers\[1\]\[49\] registers\[2\]\[49\] registers\[3\]\[49\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux4_1
XTAP_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1347 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1358 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18791_ _05045_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__buf_4
XTAP_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27989_ _12374_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1369 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_248_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_248_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17742_ registers\[4\]\[47\] registers\[5\]\[47\] registers\[6\]\[47\] registers\[7\]\[47\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__mux4_1
X_29728_ _13320_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29659_ _13284_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__clkbuf_1
X_17673_ _15830_ _04453_ _04454_ _15833_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__a22o_1
XFILLER_236_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19412_ registers\[16\]\[29\] registers\[17\]\[29\] registers\[18\]\[29\] registers\[19\]\[29\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__mux4_1
X_16624_ _15122_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
X_32670_ clknet_leaf_38_CLK _00784_ VGND VGND VPWR VPWR registers\[57\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31621_ _14316_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__clkbuf_1
X_19343_ registers\[20\]\[27\] registers\[21\]\[27\] registers\[22\]\[27\] registers\[23\]\[27\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16555_ _14952_ _15054_ _15055_ _14957_ VGND VGND VPWR VPWR _15056_ sky130_fd_sc_hd__a22o_1
XFILLER_241_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_420_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_420_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34340_ clknet_leaf_471_CLK _02454_ VGND VGND VPWR VPWR registers\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_31552_ _14280_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__clkbuf_1
X_19274_ _05844_ _06010_ _06011_ _05849_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a22o_1
X_16486_ _14985_ _14988_ _14959_ VGND VGND VPWR VPWR _14989_ sky130_fd_sc_hd__o21ba_1
XFILLER_188_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18225_ registers\[60\]\[62\] registers\[61\]\[62\] registers\[62\]\[62\] registers\[63\]\[62\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__mux4_1
X_30503_ _13728_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34271_ clknet_leaf_16_CLK _02385_ VGND VGND VPWR VPWR registers\[32\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_248_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31483_ _09762_ registers\[6\]\[34\] _14239_ VGND VGND VPWR VPWR _14244_ sky130_fd_sc_hd__mux2_1
X_36010_ clknet_leaf_407_CLK _04124_ VGND VGND VPWR VPWR registers\[63\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33222_ clknet_leaf_210_CLK _01336_ VGND VGND VPWR VPWR registers\[4\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_18156_ registers\[32\]\[60\] registers\[33\]\[60\] registers\[34\]\[60\] registers\[35\]\[60\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__mux4_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30434_ _09795_ registers\[14\]\[49\] _13682_ VGND VGND VPWR VPWR _13692_ sky130_fd_sc_hd__mux2_1
XFILLER_191_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17107_ registers\[12\]\[29\] registers\[13\]\[29\] registers\[14\]\[29\] registers\[15\]\[29\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15592_ sky130_fd_sc_hd__mux4_1
X_33153_ clknet_leaf_267_CLK _01267_ VGND VGND VPWR VPWR registers\[50\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_18087_ registers\[16\]\[57\] registers\[17\]\[57\] registers\[18\]\[57\] registers\[19\]\[57\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__mux4_2
X_30365_ _09691_ registers\[14\]\[16\] _13649_ VGND VGND VPWR VPWR _13656_ sky130_fd_sc_hd__mux2_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32104_ clknet_leaf_483_CLK _00018_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dfxtp_1
X_17038_ _15521_ _15524_ _15288_ VGND VGND VPWR VPWR _15525_ sky130_fd_sc_hd__o21ba_1
X_33084_ clknet_leaf_283_CLK _01198_ VGND VGND VPWR VPWR registers\[51\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_30296_ registers\[15\]\[48\] _13035_ _13610_ VGND VGND VPWR VPWR _13619_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_487_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_487_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_217_1244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32035_ clknet_leaf_445_CLK _00213_ VGND VGND VPWR VPWR registers\[62\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_46__f_CLK clknet_5_23_0_CLK VGND VGND VPWR VPWR clknet_6_46__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_976 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18989_ registers\[28\]\[17\] registers\[29\]\[17\] registers\[30\]\[17\] registers\[31\]\[17\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__mux4_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_239_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_239_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33986_ clknet_leaf_254_CLK _02100_ VGND VGND VPWR VPWR registers\[37\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35725_ clknet_leaf_146_CLK _03839_ VGND VGND VPWR VPWR registers\[10\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20951_ registers\[56\]\[8\] registers\[57\]\[8\] registers\[58\]\[8\] registers\[59\]\[8\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__mux4_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32937_ clknet_leaf_407_CLK _01051_ VGND VGND VPWR VPWR registers\[53\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23670_ registers\[61\]\[50\] _09797_ _09998_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__mux2_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35656_ clknet_leaf_155_CLK _03770_ VGND VGND VPWR VPWR registers\[11\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_20882_ registers\[60\]\[6\] registers\[61\]\[6\] registers\[62\]\[6\] registers\[63\]\[6\]
+ _07512_ _07329_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__mux4_1
XFILLER_148_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32868_ clknet_leaf_442_CLK _00982_ VGND VGND VPWR VPWR registers\[54\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22621_ _08953_ _09263_ _09264_ _08956_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__a22o_1
XFILLER_179_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31819_ _09660_ registers\[49\]\[1\] _14419_ VGND VGND VPWR VPWR _14421_ sky130_fd_sc_hd__mux2_1
X_34607_ clknet_leaf_411_CLK _02721_ VGND VGND VPWR VPWR registers\[27\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35587_ clknet_leaf_239_CLK _03701_ VGND VGND VPWR VPWR registers\[12\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32799_ clknet_leaf_45_CLK _00913_ VGND VGND VPWR VPWR registers\[55\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_411_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_411_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25340_ _10944_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22552_ _09194_ _09197_ _09091_ _09092_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__o211a_1
X_34538_ clknet_leaf_404_CLK _02652_ VGND VGND VPWR VPWR registers\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21503_ registers\[24\]\[23\] registers\[25\]\[23\] registers\[26\]\[23\] registers\[27\]\[23\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__mux4_1
XFILLER_194_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25271_ _10907_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__clkbuf_1
X_22483_ _09020_ _09129_ _09130_ _09024_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__a22o_1
X_34469_ clknet_leaf_464_CLK _02583_ VGND VGND VPWR VPWR registers\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_27010_ _11856_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_1
X_24222_ _09626_ registers\[58\]\[53\] _10288_ VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36208_ clknet_leaf_100_CLK _00091_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dfxtp_1
X_21434_ registers\[16\]\[21\] registers\[17\]\[21\] registers\[18\]\[21\] registers\[19\]\[21\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__mux4_1
XFILLER_124_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24153_ _09556_ registers\[58\]\[20\] _10255_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__mux2_1
X_36139_ clknet_leaf_425_CLK _04253_ VGND VGND VPWR VPWR registers\[49\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21365_ _08023_ _08030_ _08037_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__or4_2
XFILLER_200_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23104_ _09669_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20316_ registers\[52\]\[55\] registers\[53\]\[55\] registers\[54\]\[55\] registers\[55\]\[55\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__mux4_1
XFILLER_135_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24084_ _09624_ registers\[5\]\[52\] _10216_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__mux2_1
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28961_ registers\[24\]\[22\] _10351_ _12883_ VGND VGND VPWR VPWR _12886_ sky130_fd_sc_hd__mux2_1
XFILLER_174_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21296_ registers\[32\]\[18\] registers\[33\]\[18\] registers\[34\]\[18\] registers\[35\]\[18\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_478_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_478_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23035_ _09514_ VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__buf_4
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27912_ registers\[32\]\[37\] _10382_ _12326_ VGND VGND VPWR VPWR _12334_ sky130_fd_sc_hd__mux2_1
X_20247_ registers\[48\]\[53\] registers\[49\]\[53\] registers\[50\]\[53\] registers\[51\]\[53\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__mux4_1
XFILLER_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28892_ _12849_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27843_ registers\[32\]\[4\] _10313_ _12293_ VGND VGND VPWR VPWR _12298_ sky130_fd_sc_hd__mux2_1
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20178_ registers\[56\]\[51\] registers\[57\]\[51\] registers\[58\]\[51\] registers\[59\]\[51\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__mux4_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27774_ _12261_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24986_ _10726_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29513_ _09821_ registers\[21\]\[61\] _13139_ VGND VGND VPWR VPWR _13207_ sky130_fd_sc_hd__mux2_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26725_ registers\[40\]\[18\] _10342_ _11669_ VGND VGND VPWR VPWR _11678_ sky130_fd_sc_hd__mux2_1
X_23937_ _09613_ registers\[60\]\[47\] _10133_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__mux2_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_701 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_712 _07303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29444_ _09749_ registers\[21\]\[28\] _13162_ VGND VGND VPWR VPWR _13171_ sky130_fd_sc_hd__mux2_1
XFILLER_45_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_723 _07344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26656_ _11585_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__buf_4
XFILLER_166_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_734 _07356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23868_ _09544_ registers\[60\]\[14\] _10100_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__mux2_1
XANTENNA_745 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_244_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25607_ _11088_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_756 _07388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29375_ _13134_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__clkbuf_1
X_22819_ registers\[36\]\[62\] registers\[37\]\[62\] registers\[38\]\[62\] registers\[39\]\[62\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__mux4_1
XANTENNA_767 _07654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_778 _08250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26587_ _10766_ registers\[41\]\[17\] _11597_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__mux2_1
X_23799_ _09611_ registers\[29\]\[46\] _10061_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__mux2_1
XANTENNA_789 _08872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_402_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_402_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16340_ _14825_ _14832_ _14839_ _14846_ VGND VGND VPWR VPWR _14847_ sky130_fd_sc_hd__or4_4
X_28326_ registers\[2\]\[41\] _10391_ _12550_ VGND VGND VPWR VPWR _12552_ sky130_fd_sc_hd__mux2_1
X_25538_ _11050_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16271_ _14779_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__buf_2
X_28257_ _12515_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25469_ _11014_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18010_ _04683_ _04780_ _04781_ _04686_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_185_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27208_ _11780_ registers\[37\]\[24\] _11958_ VGND VGND VPWR VPWR _11963_ sky130_fd_sc_hd__mux2_1
XFILLER_139_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28188_ _12434_ VGND VGND VPWR VPWR _12479_ sky130_fd_sc_hd__buf_4
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27139_ _11926_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19961_ _06433_ _06677_ _06678_ _06439_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a22o_1
X_30150_ _13542_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18912_ registers\[12\]\[15\] registers\[13\]\[15\] registers\[14\]\[15\] registers\[15\]\[15\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_469_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_469_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19892_ _06608_ _06611_ _06504_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1100 _14530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30081_ _13494_ VGND VGND VPWR VPWR _13506_ sky130_fd_sc_hd__buf_4
XTAP_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1111 _14564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1122 _14578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18843_ _05345_ _05591_ _05592_ _05348_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__a22o_1
XANTENNA_1133 _14607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1144 _15212_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1155 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1166 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33840_ clknet_leaf_377_CLK _01954_ VGND VGND VPWR VPWR registers\[3\]\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1177 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18774_ registers\[0\]\[11\] registers\[1\]\[11\] registers\[2\]\[11\] registers\[3\]\[11\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__mux4_1
XANTENNA_1188 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _14499_ VGND VGND VPWR VPWR _14500_ sky130_fd_sc_hd__buf_12
XANTENNA_1199 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ registers\[44\]\[47\] registers\[45\]\[47\] registers\[46\]\[47\] registers\[47\]\[47\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__mux4_1
X_33771_ clknet_leaf_427_CLK _01885_ VGND VGND VPWR VPWR registers\[40\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_30983_ registers\[10\]\[53\] _13046_ _13977_ VGND VGND VPWR VPWR _13981_ sky130_fd_sc_hd__mux2_1
XFILLER_209_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32722_ clknet_leaf_174_CLK _00836_ VGND VGND VPWR VPWR registers\[56\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35510_ clknet_leaf_319_CLK _03624_ VGND VGND VPWR VPWR registers\[13\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17656_ registers\[36\]\[45\] registers\[37\]\[45\] registers\[38\]\[45\] registers\[39\]\[45\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__mux4_1
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16607_ _14502_ VGND VGND VPWR VPWR _15106_ sky130_fd_sc_hd__buf_4
X_35441_ clknet_leaf_377_CLK _03555_ VGND VGND VPWR VPWR registers\[14\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32653_ clknet_leaf_139_CLK _00767_ VGND VGND VPWR VPWR registers\[58\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17587_ registers\[32\]\[43\] registers\[33\]\[43\] registers\[34\]\[43\] registers\[35\]\[43\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__mux4_1
XFILLER_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31604_ _14307_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__clkbuf_1
X_19326_ registers\[48\]\[27\] registers\[49\]\[27\] registers\[50\]\[27\] registers\[51\]\[27\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__mux4_1
X_16538_ registers\[52\]\[13\] registers\[53\]\[13\] registers\[54\]\[13\] registers\[55\]\[13\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _15039_ sky130_fd_sc_hd__mux4_1
X_35372_ clknet_leaf_394_CLK _03486_ VGND VGND VPWR VPWR registers\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32584_ clknet_leaf_160_CLK _00698_ VGND VGND VPWR VPWR registers\[5\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34323_ clknet_leaf_103_CLK _02437_ VGND VGND VPWR VPWR registers\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_31535_ _09817_ registers\[6\]\[59\] _14261_ VGND VGND VPWR VPWR _14271_ sky130_fd_sc_hd__mux2_1
XFILLER_148_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19257_ registers\[52\]\[25\] registers\[53\]\[25\] registers\[54\]\[25\] registers\[55\]\[25\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__mux4_1
X_16469_ registers\[60\]\[11\] registers\[61\]\[11\] registers\[62\]\[11\] registers\[63\]\[11\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _14972_ sky130_fd_sc_hd__mux4_1
XFILLER_223_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18208_ _14558_ _04972_ _04973_ _14568_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__a22o_1
X_34254_ clknet_leaf_131_CLK _02368_ VGND VGND VPWR VPWR registers\[32\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31466_ _09744_ registers\[6\]\[26\] _14228_ VGND VGND VPWR VPWR _14235_ sky130_fd_sc_hd__mux2_1
X_19188_ registers\[48\]\[23\] registers\[49\]\[23\] registers\[50\]\[23\] registers\[51\]\[23\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__mux4_1
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33205_ clknet_leaf_321_CLK _01319_ VGND VGND VPWR VPWR registers\[4\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_18139_ registers\[8\]\[59\] registers\[9\]\[59\] registers\[10\]\[59\] registers\[11\]\[59\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30417_ _13683_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__clkbuf_1
X_34185_ clknet_leaf_238_CLK _02299_ VGND VGND VPWR VPWR registers\[34\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_31397_ _14198_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33136_ clknet_leaf_366_CLK _01250_ VGND VGND VPWR VPWR registers\[50\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_21150_ registers\[24\]\[13\] registers\[25\]\[13\] registers\[26\]\[13\] registers\[27\]\[13\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__mux4_1
XFILLER_171_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30348_ _09674_ registers\[14\]\[8\] _13638_ VGND VGND VPWR VPWR _13647_ sky130_fd_sc_hd__mux2_1
X_20101_ _06576_ _06813_ _06814_ _06579_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__a22o_1
XFILLER_67_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21081_ registers\[16\]\[11\] registers\[17\]\[11\] registers\[18\]\[11\] registers\[19\]\[11\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__mux4_1
X_33067_ clknet_leaf_419_CLK _01181_ VGND VGND VPWR VPWR registers\[51\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30279_ _13565_ VGND VGND VPWR VPWR _13610_ sky130_fd_sc_hd__buf_4
XFILLER_193_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32018_ clknet_leaf_64_CLK _00196_ VGND VGND VPWR VPWR registers\[62\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_20032_ registers\[48\]\[47\] registers\[49\]\[47\] registers\[50\]\[47\] registers\[51\]\[47\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__mux4_1
XFILLER_140_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24840_ _09634_ registers\[54\]\[57\] _10642_ VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__mux2_1
XFILLER_86_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21983_ _08334_ _08643_ _08644_ _08338_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__a22o_1
X_24771_ _09565_ registers\[54\]\[24\] _10609_ VGND VGND VPWR VPWR _10614_ sky130_fd_sc_hd__mux2_1
XFILLER_67_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33969_ clknet_leaf_358_CLK _02083_ VGND VGND VPWR VPWR registers\[37\]\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26510_ _10825_ registers\[42\]\[45\] _11558_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__mux2_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35708_ clknet_leaf_300_CLK _03822_ VGND VGND VPWR VPWR registers\[10\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_23722_ _10027_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
X_20934_ registers\[16\]\[7\] registers\[17\]\[7\] registers\[18\]\[7\] registers\[19\]\[7\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__mux4_1
XFILLER_27_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27490_ _12077_ VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__buf_4
XFILLER_187_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26441_ _10756_ registers\[42\]\[12\] _11525_ VGND VGND VPWR VPWR _11528_ sky130_fd_sc_hd__mux2_1
X_20865_ _07373_ _07557_ _07558_ _07383_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__a22o_1
X_23653_ registers\[61\]\[42\] _09780_ _09987_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__mux2_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35639_ clknet_leaf_318_CLK _03753_ VGND VGND VPWR VPWR registers\[11\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_880 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22604_ _09248_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29160_ net29 VGND VGND VPWR VPWR _13008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23584_ _09953_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
X_26372_ _11491_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__clkbuf_1
X_20796_ _07486_ _07491_ _07370_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__o21ba_1
XFILLER_165_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28111_ _11736_ registers\[30\]\[3\] _12435_ VGND VGND VPWR VPWR _12439_ sky130_fd_sc_hd__mux2_1
XFILLER_10_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22535_ _09109_ _09180_ _09181_ _09114_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__a22o_1
X_25323_ _10934_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29091_ _12961_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28042_ _12402_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__clkbuf_1
X_22466_ _09109_ _09110_ _09113_ _09114_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__a22o_1
XFILLER_182_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25254_ _10793_ registers\[51\]\[30\] _10898_ VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__mux2_1
XFILLER_136_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24205_ _09609_ registers\[58\]\[45\] _10277_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__mux2_1
X_21417_ _07783_ _08093_ _08094_ _07786_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__a22o_1
X_25185_ _10861_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__clkbuf_1
X_22397_ registers\[32\]\[49\] registers\[33\]\[49\] registers\[34\]\[49\] registers\[35\]\[49\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__mux4_1
XFILLER_68_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24136_ _09540_ registers\[58\]\[12\] _10244_ VGND VGND VPWR VPWR _10247_ sky130_fd_sc_hd__mux2_1
XFILLER_120_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21348_ registers\[52\]\[19\] registers\[53\]\[19\] registers\[54\]\[19\] registers\[55\]\[19\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__mux4_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29993_ registers\[17\]\[32\] _13002_ _13457_ VGND VGND VPWR VPWR _13460_ sky130_fd_sc_hd__mux2_1
XFILLER_151_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24067_ _09607_ registers\[5\]\[44\] _10205_ VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__mux2_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28944_ registers\[24\]\[14\] _10334_ _12872_ VGND VGND VPWR VPWR _12877_ sky130_fd_sc_hd__mux2_1
X_21279_ registers\[8\]\[17\] registers\[9\]\[17\] registers\[10\]\[17\] registers\[11\]\[17\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23018_ _09608_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28875_ _12840_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27826_ _12288_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__clkbuf_1
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27757_ _12252_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__clkbuf_1
X_24969_ _09628_ registers\[53\]\[54\] _10713_ VGND VGND VPWR VPWR _10718_ sky130_fd_sc_hd__mux2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17510_ _14544_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__clkbuf_4
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26708_ _11657_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__buf_4
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18490_ _05107_ _05248_ _05249_ _05117_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__a22o_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27688_ registers\[34\]\[59\] _10428_ _12206_ VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__mux2_1
XFILLER_206_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_520 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_531 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_542 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29427_ _13139_ VGND VGND VPWR VPWR _13162_ sky130_fd_sc_hd__buf_4
XFILLER_79_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17441_ registers\[40\]\[39\] registers\[41\]\[39\] registers\[42\]\[39\] registers\[43\]\[39\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15916_ sky130_fd_sc_hd__mux4_1
XFILLER_221_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_553 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26639_ _11632_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_564 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_575 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_586 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29358_ _09800_ registers\[22\]\[51\] _13124_ VGND VGND VPWR VPWR _13126_ sky130_fd_sc_hd__mux2_1
XANTENNA_597 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17372_ registers\[44\]\[37\] registers\[45\]\[37\] registers\[46\]\[37\] registers\[47\]\[37\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15849_ sky130_fd_sc_hd__mux4_1
XFILLER_92_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19111_ _05853_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16323_ registers\[52\]\[7\] registers\[53\]\[7\] registers\[54\]\[7\] registers\[55\]\[7\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14830_ sky130_fd_sc_hd__mux4_1
X_28309_ registers\[2\]\[33\] _10374_ _12539_ VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__mux2_1
XFILLER_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29289_ _13089_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31320_ _14158_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19042_ _05547_ _05784_ _05785_ _05550_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a22o_1
XFILLER_174_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16254_ _14502_ VGND VGND VPWR VPWR _14763_ sky130_fd_sc_hd__buf_6
XFILLER_71_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31251_ registers\[8\]\[52\] net48 _14119_ VGND VGND VPWR VPWR _14122_ sky130_fd_sc_hd__mux2_1
XFILLER_138_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16185_ registers\[52\]\[3\] registers\[53\]\[3\] registers\[54\]\[3\] registers\[55\]\[3\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14696_ sky130_fd_sc_hd__mux4_1
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 net207 VGND VGND VPWR VPWR D2[58] sky130_fd_sc_hd__buf_2
X_30202_ registers\[15\]\[3\] _12941_ _13566_ VGND VGND VPWR VPWR _13570_ sky130_fd_sc_hd__mux2_1
Xoutput218 net218 VGND VGND VPWR VPWR D3[0] sky130_fd_sc_hd__buf_2
XFILLER_138_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31182_ _14085_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__clkbuf_1
Xoutput229 net229 VGND VGND VPWR VPWR D3[1] sky130_fd_sc_hd__buf_2
XFILLER_245_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30133_ _13533_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19944_ registers\[16\]\[44\] registers\[17\]\[44\] registers\[18\]\[44\] registers\[19\]\[44\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__mux4_1
X_35990_ clknet_leaf_184_CLK _04104_ VGND VGND VPWR VPWR registers\[63\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30064_ _13497_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__clkbuf_1
X_34941_ clknet_leaf_186_CLK _03055_ VGND VGND VPWR VPWR registers\[22\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_19875_ registers\[24\]\[42\] registers\[25\]\[42\] registers\[26\]\[42\] registers\[27\]\[42\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__mux4_1
XFILLER_150_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18826_ _05576_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
XTAP_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34872_ clknet_leaf_309_CLK _02986_ VGND VGND VPWR VPWR registers\[23\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33823_ clknet_leaf_486_CLK _01937_ VGND VGND VPWR VPWR registers\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_18757_ _05476_ _05485_ _05495_ _05509_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__or4_2
XFILLER_236_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17708_ _14581_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__buf_4
XFILLER_97_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33754_ clknet_leaf_32_CLK _01868_ VGND VGND VPWR VPWR registers\[40\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_18688_ registers\[36\]\[9\] registers\[37\]\[9\] registers\[38\]\[9\] registers\[39\]\[9\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__mux4_1
X_30966_ registers\[10\]\[45\] _13029_ _13966_ VGND VGND VPWR VPWR _13972_ sky130_fd_sc_hd__mux2_1
XFILLER_110_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32705_ clknet_leaf_266_CLK _00819_ VGND VGND VPWR VPWR registers\[57\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17639_ _15830_ _04420_ _04421_ _15833_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__a22o_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33685_ clknet_leaf_125_CLK _01799_ VGND VGND VPWR VPWR registers\[41\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30897_ registers\[10\]\[12\] _12960_ _13933_ VGND VGND VPWR VPWR _13936_ sky130_fd_sc_hd__mux2_1
XFILLER_212_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32636_ clknet_leaf_289_CLK _00750_ VGND VGND VPWR VPWR registers\[58\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_20650_ _07316_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__buf_12
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35424_ clknet_leaf_483_CLK _03538_ VGND VGND VPWR VPWR registers\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19309_ _05839_ _06042_ _06045_ _05842_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__a22o_1
XFILLER_177_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35355_ clknet_leaf_477_CLK _03469_ VGND VGND VPWR VPWR registers\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_20581_ net72 VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__buf_8
XFILLER_220_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32567_ clknet_leaf_313_CLK _00681_ VGND VGND VPWR VPWR registers\[5\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22320_ _08943_ _08952_ _08963_ _08972_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__or4_4
XFILLER_104_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34306_ clknet_leaf_249_CLK _02420_ VGND VGND VPWR VPWR registers\[32\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_31518_ _14262_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35286_ clknet_leaf_86_CLK _03400_ VGND VGND VPWR VPWR registers\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32498_ clknet_leaf_379_CLK _00612_ VGND VGND VPWR VPWR registers\[60\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34237_ clknet_leaf_278_CLK _02351_ VGND VGND VPWR VPWR registers\[33\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_22251_ _08905_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_2
XFILLER_192_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31449_ _09695_ registers\[6\]\[18\] _14217_ VGND VGND VPWR VPWR _14226_ sky130_fd_sc_hd__mux2_1
XFILLER_191_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21202_ _07640_ _07884_ _07885_ _07646_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__a22o_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22182_ _08766_ _08837_ _08838_ _08771_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__a22o_1
X_34168_ clknet_leaf_337_CLK _02282_ VGND VGND VPWR VPWR registers\[34\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33119_ clknet_leaf_36_CLK _01233_ VGND VGND VPWR VPWR registers\[50\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_21133_ _07815_ _07818_ _07711_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__o21ba_1
XFILLER_156_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26990_ net50 VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__buf_4
X_34099_ clknet_leaf_349_CLK _02213_ VGND VGND VPWR VPWR registers\[35\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21064_ _07440_ _07750_ _07751_ _07443_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a22o_1
X_25941_ _10796_ registers\[46\]\[31\] _11263_ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__mux2_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20015_ _06525_ _06728_ _06731_ _06528_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__a22o_1
XFILLER_154_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28660_ _12727_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25872_ _10862_ registers\[47\]\[63\] _11158_ VGND VGND VPWR VPWR _11228_ sky130_fd_sc_hd__mux2_1
XFILLER_87_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27611_ registers\[34\]\[22\] _10351_ _12173_ VGND VGND VPWR VPWR _12176_ sky130_fd_sc_hd__mux2_1
X_24823_ _09617_ registers\[54\]\[49\] _10631_ VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28591_ _11811_ registers\[27\]\[39\] _12681_ VGND VGND VPWR VPWR _12691_ sky130_fd_sc_hd__mux2_1
XFILLER_246_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27542_ _12138_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__clkbuf_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24754_ _09548_ registers\[54\]\[16\] _10598_ VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__mux2_1
X_21966_ _08625_ _08628_ _08430_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__o21ba_1
XFILLER_243_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23705_ _09517_ registers\[29\]\[1\] _10017_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__mux2_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20917_ _07440_ _07605_ _07608_ _07443_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__a22o_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27473_ _12102_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24685_ _10567_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
X_21897_ _08536_ _08545_ _08552_ _08561_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__or4_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29212_ _13043_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26424_ _10739_ registers\[42\]\[4\] _11514_ VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__mux2_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20848_ registers\[48\]\[5\] registers\[49\]\[5\] registers\[50\]\[5\] registers\[51\]\[5\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__mux4_1
X_23636_ registers\[61\]\[34\] _09762_ _09976_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__mux2_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29143_ _12996_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26355_ _11482_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__clkbuf_1
X_20779_ _07440_ _07473_ _07474_ _07443_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__a22o_1
X_23567_ registers\[61\]\[1\] _09660_ _09943_ VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25306_ _10846_ registers\[51\]\[55\] _10920_ VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__mux2_1
X_22518_ registers\[52\]\[52\] registers\[53\]\[52\] registers\[54\]\[52\] registers\[55\]\[52\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__mux4_1
X_29074_ registers\[23\]\[7\] _12949_ _12935_ VGND VGND VPWR VPWR _12950_ sky130_fd_sc_hd__mux2_1
X_26286_ _11446_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
X_23498_ _09907_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28025_ _12393_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__clkbuf_1
X_22449_ _08953_ _09094_ _09097_ _08956_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__a22o_1
XFILLER_13_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25237_ _10777_ registers\[51\]\[22\] _10887_ VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__mux2_1
XFILLER_183_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25168_ net53 VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__buf_4
XFILLER_164_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24119_ _09523_ registers\[58\]\[4\] _10233_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__mux2_1
XFILLER_150_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17990_ registers\[12\]\[54\] registers\[13\]\[54\] registers\[14\]\[54\] registers\[15\]\[54\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__mux4_1
X_25099_ _10803_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__clkbuf_1
X_29976_ registers\[17\]\[24\] _12985_ _13446_ VGND VGND VPWR VPWR _13451_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28927_ registers\[24\]\[6\] _10317_ _12861_ VGND VGND VPWR VPWR _12868_ sky130_fd_sc_hd__mux2_1
X_16941_ registers\[20\]\[24\] registers\[21\]\[24\] registers\[22\]\[24\] registers\[23\]\[24\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15431_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19660_ _05081_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__buf_4
XFILLER_77_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16872_ _14592_ VGND VGND VPWR VPWR _15364_ sky130_fd_sc_hd__buf_4
X_28858_ _12831_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18611_ registers\[32\]\[7\] registers\[33\]\[7\] registers\[34\]\[7\] registers\[35\]\[7\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__mux4_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27809_ registers\[33\]\[52\] _10414_ _12277_ VGND VGND VPWR VPWR _12280_ sky130_fd_sc_hd__mux2_1
XFILLER_219_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19591_ registers\[16\]\[34\] registers\[17\]\[34\] registers\[18\]\[34\] registers\[19\]\[34\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__mux4_1
XFILLER_231_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28789_ _12795_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__clkbuf_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _05197_ _05298_ _05299_ _05202_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a22o_1
X_30820_ _13850_ VGND VGND VPWR VPWR _13895_ sky130_fd_sc_hd__buf_4
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30751_ _09672_ registers\[11\]\[7\] _13851_ VGND VGND VPWR VPWR _13859_ sky130_fd_sc_hd__mux2_1
X_18473_ _05233_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__clkbuf_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_372 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17424_ registers\[0\]\[38\] registers\[1\]\[38\] registers\[2\]\[38\] registers\[3\]\[38\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15900_ sky130_fd_sc_hd__mux4_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33470_ clknet_leaf_273_CLK _01584_ VGND VGND VPWR VPWR registers\[45\]\[48\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_383 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30682_ _13822_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_394 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32421_ clknet_leaf_464_CLK _00535_ VGND VGND VPWR VPWR registers\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _14581_ VGND VGND VPWR VPWR _15833_ sky130_fd_sc_hd__buf_4
XFILLER_140_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35140_ clknet_leaf_224_CLK _03254_ VGND VGND VPWR VPWR registers\[1\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16306_ _14601_ _14812_ _14813_ _14611_ VGND VGND VPWR VPWR _14814_ sky130_fd_sc_hd__a22o_1
X_32352_ clknet_leaf_44_CLK _00466_ VGND VGND VPWR VPWR registers\[61\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_17286_ _15487_ _15764_ _15765_ _15490_ VGND VGND VPWR VPWR _15766_ sky130_fd_sc_hd__a22o_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19025_ _05764_ _05769_ _05494_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__o21ba_1
X_31303_ _14149_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16237_ _14743_ _14746_ _14614_ VGND VGND VPWR VPWR _14747_ sky130_fd_sc_hd__o21ba_1
X_35071_ clknet_leaf_305_CLK _03185_ VGND VGND VPWR VPWR registers\[20\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_32283_ clknet_leaf_20_CLK _00397_ VGND VGND VPWR VPWR registers\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34022_ clknet_leaf_434_CLK _02136_ VGND VGND VPWR VPWR registers\[36\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31234_ registers\[8\]\[44\] net39 _14108_ VGND VGND VPWR VPWR _14113_ sky130_fd_sc_hd__mux2_1
X_16168_ registers\[28\]\[2\] registers\[29\]\[2\] registers\[30\]\[2\] registers\[31\]\[2\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14680_ sky130_fd_sc_hd__mux4_1
XFILLER_127_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31165_ registers\[8\]\[11\] net3 _14075_ VGND VGND VPWR VPWR _14077_ sky130_fd_sc_hd__mux2_1
X_16099_ net70 net69 VGND VGND VPWR VPWR _14613_ sky130_fd_sc_hd__or2b_4
XFILLER_173_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30116_ _13524_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19927_ registers\[48\]\[44\] registers\[49\]\[44\] registers\[50\]\[44\] registers\[51\]\[44\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__mux4_1
XFILLER_229_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35973_ clknet_leaf_230_CLK _04087_ VGND VGND VPWR VPWR registers\[6\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31096_ _14040_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30047_ registers\[17\]\[58\] _13056_ _13479_ VGND VGND VPWR VPWR _13488_ sky130_fd_sc_hd__mux2_1
X_34924_ clknet_leaf_402_CLK _03038_ VGND VGND VPWR VPWR registers\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19858_ _05065_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_151_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18809_ registers\[8\]\[12\] registers\[9\]\[12\] registers\[10\]\[12\] registers\[11\]\[12\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__mux4_1
X_34855_ clknet_leaf_455_CLK _02969_ VGND VGND VPWR VPWR registers\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_216_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19789_ _05102_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33806_ clknet_leaf_109_CLK _01920_ VGND VGND VPWR VPWR registers\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_21820_ _08272_ _08485_ _08486_ _08275_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__a22o_1
XFILLER_3_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31998_ clknet_leaf_29_CLK _00170_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_1
X_34786_ clknet_leaf_446_CLK _02900_ VGND VGND VPWR VPWR registers\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21751_ registers\[16\]\[30\] registers\[17\]\[30\] registers\[18\]\[30\] registers\[19\]\[30\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__mux4_1
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33737_ clknet_leaf_245_CLK _01851_ VGND VGND VPWR VPWR registers\[41\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30949_ registers\[10\]\[37\] _13012_ _13955_ VGND VGND VPWR VPWR _13963_ sky130_fd_sc_hd__mux2_1
XFILLER_52_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20702_ _07311_ _07342_ _07371_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__or4_4
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24470_ _10453_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
X_21682_ registers\[28\]\[28\] registers\[29\]\[28\] registers\[30\]\[28\] registers\[31\]\[28\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__mux4_1
X_33668_ clknet_leaf_251_CLK _01782_ VGND VGND VPWR VPWR registers\[42\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35407_ clknet_leaf_137_CLK _03521_ VGND VGND VPWR VPWR registers\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_23421_ registers\[39\]\[63\] _09825_ _09657_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__mux2_1
X_20633_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__buf_4
XFILLER_36_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32619_ clknet_leaf_420_CLK _00733_ VGND VGND VPWR VPWR registers\[58\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_33599_ clknet_leaf_272_CLK _01713_ VGND VGND VPWR VPWR registers\[43\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26140_ _10860_ registers\[45\]\[62\] _11300_ VGND VGND VPWR VPWR _11369_ sky130_fd_sc_hd__mux2_1
XFILLER_177_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23352_ _09657_ VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__buf_4
X_35338_ clknet_leaf_149_CLK _03452_ VGND VGND VPWR VPWR registers\[16\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_20564_ _05060_ _07262_ _07263_ _05066_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__a22o_1
XFILLER_221_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22303_ _07352_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__buf_4
XFILLER_165_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23283_ net39 VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__clkbuf_4
X_26071_ _10791_ registers\[45\]\[29\] _11323_ VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__mux2_1
X_35269_ clknet_leaf_220_CLK _03383_ VGND VGND VPWR VPWR registers\[17\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_20495_ registers\[60\]\[61\] registers\[61\]\[61\] registers\[62\]\[61\] registers\[63\]\[61\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__mux4_1
XFILLER_192_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_23_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_23_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22234_ registers\[8\]\[44\] registers\[9\]\[44\] registers\[10\]\[44\] registers\[11\]\[44\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__mux4_1
X_25022_ net2 VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__buf_2
XFILLER_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29830_ registers\[18\]\[19\] _12974_ _13364_ VGND VGND VPWR VPWR _13374_ sky130_fd_sc_hd__mux2_1
X_22165_ registers\[52\]\[42\] registers\[53\]\[42\] registers\[54\]\[42\] registers\[55\]\[42\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__mux4_1
XTAP_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21116_ registers\[24\]\[12\] registers\[25\]\[12\] registers\[26\]\[12\] registers\[27\]\[12\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__mux4_1
XTAP_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29761_ registers\[1\]\[50\] _13039_ _13337_ VGND VGND VPWR VPWR _13338_ sky130_fd_sc_hd__mux2_1
XFILLER_133_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26973_ _11831_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_1
X_22096_ _08610_ _08751_ _08754_ _08613_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__a22o_1
XTAP_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28712_ _11797_ registers\[26\]\[32\] _12752_ VGND VGND VPWR VPWR _12755_ sky130_fd_sc_hd__mux2_1
X_25924_ _10779_ registers\[46\]\[23\] _11252_ VGND VGND VPWR VPWR _11256_ sky130_fd_sc_hd__mux2_1
X_21047_ _07732_ _07733_ _07734_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__a22o_1
X_29692_ _13301_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28643_ _10014_ _10935_ VGND VGND VPWR VPWR _12718_ sky130_fd_sc_hd__nand2_8
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25855_ _11219_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24806_ _10632_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28574_ _12682_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__clkbuf_1
X_25786_ _11183_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
X_22998_ _09594_ registers\[62\]\[38\] _09578_ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__mux2_1
X_27525_ _12129_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__clkbuf_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ _09531_ registers\[54\]\[8\] _10587_ VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__mux2_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ registers\[0\]\[36\] registers\[1\]\[36\] registers\[2\]\[36\] registers\[3\]\[36\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__mux4_1
XFILLER_215_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27456_ _12093_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__clkbuf_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _09598_ registers\[55\]\[40\] _10558_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__mux2_1
XFILLER_199_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26407_ _11509_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__clkbuf_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23619_ registers\[61\]\[26\] _09744_ _09965_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__mux2_1
XFILLER_230_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27387_ registers\[36\]\[45\] _10399_ _12051_ VGND VGND VPWR VPWR _12057_ sky130_fd_sc_hd__mux2_1
XFILLER_129_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24599_ _10522_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_927 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29126_ net17 VGND VGND VPWR VPWR _12985_ sky130_fd_sc_hd__buf_2
X_17140_ _14562_ VGND VGND VPWR VPWR _15624_ sky130_fd_sc_hd__buf_6
X_26338_ _11473_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29057_ _12938_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17071_ registers\[0\]\[28\] registers\[1\]\[28\] registers\[2\]\[28\] registers\[3\]\[28\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15557_ sky130_fd_sc_hd__mux4_1
X_26269_ _10854_ registers\[44\]\[59\] _11427_ VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__mux2_1
XFILLER_7_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16022_ registers\[48\]\[0\] registers\[49\]\[0\] registers\[50\]\[0\] registers\[51\]\[0\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14536_ sky130_fd_sc_hd__mux4_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28008_ _12384_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17973_ _04676_ _04744_ _04745_ _04681_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a22o_1
XFILLER_151_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29959_ registers\[17\]\[16\] _12968_ _13435_ VGND VGND VPWR VPWR _13442_ sky130_fd_sc_hd__mux2_1
XFILLER_97_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16924_ registers\[60\]\[24\] registers\[61\]\[24\] registers\[62\]\[24\] registers\[63\]\[24\]
+ _15413_ _15207_ VGND VGND VPWR VPWR _15414_ sky130_fd_sc_hd__mux4_1
X_19712_ _05092_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__clkbuf_4
X_32970_ clknet_leaf_162_CLK _01084_ VGND VGND VPWR VPWR registers\[53\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31921_ _14418_ VGND VGND VPWR VPWR _14474_ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16855_ registers\[56\]\[22\] registers\[57\]\[22\] registers\[58\]\[22\] registers\[59\]\[22\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15347_ sky130_fd_sc_hd__mux4_1
X_19643_ _05097_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__buf_4
XFILLER_226_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34640_ clknet_leaf_116_CLK _02754_ VGND VGND VPWR VPWR registers\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19574_ registers\[48\]\[34\] registers\[49\]\[34\] registers\[50\]\[34\] registers\[51\]\[34\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__mux4_1
XFILLER_53_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31852_ _09693_ registers\[49\]\[17\] _14430_ VGND VGND VPWR VPWR _14438_ sky130_fd_sc_hd__mux2_1
XFILLER_225_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16786_ registers\[8\]\[20\] registers\[9\]\[20\] registers\[10\]\[20\] registers\[11\]\[20\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15280_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18525_ registers\[12\]\[4\] registers\[13\]\[4\] registers\[14\]\[4\] registers\[15\]\[4\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__mux4_1
X_30803_ _13886_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34571_ clknet_leaf_158_CLK _02685_ VGND VGND VPWR VPWR registers\[28\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31783_ _14401_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30734_ _13849_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__clkbuf_1
X_18456_ registers\[8\]\[2\] registers\[9\]\[2\] registers\[10\]\[2\] registers\[11\]\[2\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux4_1
X_33522_ clknet_leaf_361_CLK _01636_ VGND VGND VPWR VPWR registers\[44\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_180 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_191 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17407_ _15879_ _15882_ _15612_ VGND VGND VPWR VPWR _15883_ sky130_fd_sc_hd__o21ba_1
X_33453_ clknet_leaf_345_CLK _01567_ VGND VGND VPWR VPWR registers\[45\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_18387_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__buf_4
X_30665_ registers\[12\]\[30\] _12997_ _13813_ VGND VGND VPWR VPWR _13814_ sky130_fd_sc_hd__mux2_1
XFILLER_226_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32404_ clknet_leaf_93_CLK _00518_ VGND VGND VPWR VPWR registers\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17338_ registers\[56\]\[36\] registers\[57\]\[36\] registers\[58\]\[36\] registers\[59\]\[36\]
+ _15752_ _15542_ VGND VGND VPWR VPWR _15816_ sky130_fd_sc_hd__mux4_1
X_36172_ clknet_leaf_168_CLK _04286_ VGND VGND VPWR VPWR registers\[49\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33384_ clknet_leaf_59_CLK _01498_ VGND VGND VPWR VPWR registers\[46\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_30596_ _09823_ registers\[13\]\[62\] _13708_ VGND VGND VPWR VPWR _13777_ sky130_fd_sc_hd__mux2_1
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32335_ clknet_leaf_172_CLK _00449_ VGND VGND VPWR VPWR registers\[61\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_35123_ clknet_leaf_384_CLK _03237_ VGND VGND VPWR VPWR registers\[1\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17269_ registers\[36\]\[34\] registers\[37\]\[34\] registers\[38\]\[34\] registers\[39\]\[34\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15749_ sky130_fd_sc_hd__mux4_1
XFILLER_105_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19008_ _05049_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35054_ clknet_leaf_387_CLK _03168_ VGND VGND VPWR VPWR registers\[20\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_32266_ clknet_leaf_159_CLK _00380_ VGND VGND VPWR VPWR registers\[39\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_20280_ registers\[48\]\[54\] registers\[49\]\[54\] registers\[50\]\[54\] registers\[51\]\[54\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__mux4_1
XFILLER_146_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34005_ clknet_leaf_120_CLK _02119_ VGND VGND VPWR VPWR registers\[36\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_31217_ registers\[8\]\[36\] net30 _14097_ VGND VGND VPWR VPWR _14104_ sky130_fd_sc_hd__mux2_1
X_32197_ clknet_leaf_391_CLK _00311_ VGND VGND VPWR VPWR registers\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31148_ registers\[8\]\[3\] net34 _14064_ VGND VGND VPWR VPWR _14068_ sky130_fd_sc_hd__mux2_1
XFILLER_170_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23970_ _09646_ registers\[60\]\[63\] _10088_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__mux2_1
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31079_ _14031_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__clkbuf_1
X_35956_ clknet_leaf_321_CLK _04070_ VGND VGND VPWR VPWR registers\[6\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22921_ _09542_ registers\[62\]\[13\] _09536_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34907_ clknet_leaf_490_CLK _03021_ VGND VGND VPWR VPWR registers\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35887_ clknet_leaf_378_CLK _04001_ VGND VGND VPWR VPWR registers\[7\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25640_ _11105_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
X_22852_ registers\[56\]\[63\] registers\[57\]\[63\] registers\[58\]\[63\] registers\[59\]\[63\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__mux4_1
X_34838_ clknet_leaf_97_CLK _02952_ VGND VGND VPWR VPWR registers\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21803_ registers\[44\]\[32\] registers\[45\]\[32\] registers\[46\]\[32\] registers\[47\]\[32\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__mux4_1
X_25571_ registers\[4\]\[50\] _10409_ _11067_ VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__mux2_1
X_22783_ _09400_ _09407_ _09414_ _09421_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__or4_4
X_34769_ clknet_leaf_111_CLK _02883_ VGND VGND VPWR VPWR registers\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_27310_ _12016_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__clkbuf_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24522_ _10480_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28290_ registers\[2\]\[24\] _10355_ _12528_ VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__mux2_1
X_21734_ registers\[52\]\[30\] registers\[53\]\[30\] registers\[54\]\[30\] registers\[55\]\[30\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__mux4_1
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27241_ _11935_ VGND VGND VPWR VPWR _11980_ sky130_fd_sc_hd__buf_4
X_24453_ _10444_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21665_ registers\[60\]\[28\] registers\[61\]\[28\] registers\[62\]\[28\] registers\[63\]\[28\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__mux4_1
XFILLER_200_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23404_ _09856_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
X_27172_ _11744_ registers\[37\]\[7\] _11936_ VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20616_ _07314_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__buf_12
XFILLER_177_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24384_ _10398_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
X_21596_ registers\[0\]\[26\] registers\[1\]\[26\] registers\[2\]\[26\] registers\[3\]\[26\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__mux4_1
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26123_ _11360_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23335_ _09818_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
X_20547_ _05077_ _07245_ _07246_ _05086_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__a22o_1
XFILLER_197_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26054_ _11324_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
X_20478_ _05107_ _07179_ _07180_ _05117_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__a22o_1
X_23266_ _09772_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25005_ _10739_ registers\[52\]\[4\] _10731_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__mux2_1
X_22217_ _08872_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_2
X_23197_ registers\[9\]\[16\] _09691_ _09722_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__mux2_1
XFILLER_134_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22148_ _07312_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__clkbuf_4
X_29813_ _13365_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1507 _07382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1518 _08841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1529 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29744_ registers\[1\]\[42\] _13023_ _13326_ VGND VGND VPWR VPWR _13329_ sky130_fd_sc_hd__mux2_1
X_26956_ net38 VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__buf_4
X_22079_ registers\[36\]\[40\] registers\[37\]\[40\] registers\[38\]\[40\] registers\[39\]\[40\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__mux4_1
XTAP_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25907_ _10762_ registers\[46\]\[15\] _11241_ VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__mux2_1
X_29675_ _13292_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26887_ _11773_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28626_ _12709_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ _15132_ _15137_ _14934_ _14935_ VGND VGND VPWR VPWR _15138_ sky130_fd_sc_hd__o211a_2
XFILLER_247_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25838_ _11210_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28557_ _12673_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__clkbuf_1
X_16571_ registers\[60\]\[14\] registers\[61\]\[14\] registers\[62\]\[14\] registers\[63\]\[14\]
+ _15070_ _14864_ VGND VGND VPWR VPWR _15071_ sky130_fd_sc_hd__mux4_1
X_25769_ _11174_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18310_ net81 net82 VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__or2b_4
XFILLER_128_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27508_ _12120_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__clkbuf_1
X_19290_ _05097_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__buf_6
XFILLER_215_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28488_ _11843_ registers\[28\]\[54\] _12632_ VGND VGND VPWR VPWR _12637_ sky130_fd_sc_hd__mux2_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _14570_ _05004_ _05005_ _14582_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__a22o_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27439_ _12084_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18172_ registers\[12\]\[60\] registers\[13\]\[60\] registers\[14\]\[60\] registers\[15\]\[60\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__mux4_1
X_30450_ _13700_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29109_ _12973_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__clkbuf_1
X_17123_ _14546_ VGND VGND VPWR VPWR _15607_ sky130_fd_sc_hd__buf_4
XFILLER_106_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30381_ _13664_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32120_ clknet_leaf_465_CLK _00036_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17054_ _15536_ _15539_ _15269_ VGND VGND VPWR VPWR _15540_ sky130_fd_sc_hd__o21ba_1
XFILLER_7_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16005_ _14518_ VGND VGND VPWR VPWR _14519_ sky130_fd_sc_hd__buf_4
X_32051_ clknet_leaf_379_CLK _00229_ VGND VGND VPWR VPWR registers\[62\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31002_ _13990_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__clkbuf_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35810_ clknet_leaf_465_CLK _03924_ VGND VGND VPWR VPWR registers\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17956_ _14518_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__buf_6
XFILLER_112_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35741_ clknet_leaf_478_CLK _03855_ VGND VGND VPWR VPWR registers\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_16907_ registers\[20\]\[23\] registers\[21\]\[23\] registers\[22\]\[23\] registers\[23\]\[23\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15398_ sky130_fd_sc_hd__mux4_1
X_17887_ _04481_ _04661_ _04662_ _04484_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a22o_1
X_32953_ clknet_leaf_286_CLK _01067_ VGND VGND VPWR VPWR registers\[53\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19626_ registers\[20\]\[35\] registers\[21\]\[35\] registers\[22\]\[35\] registers\[23\]\[35\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__mux4_1
X_31904_ _14465_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__clkbuf_1
X_16838_ _15295_ _15329_ _15330_ _15300_ VGND VGND VPWR VPWR _15331_ sky130_fd_sc_hd__a22o_1
X_35672_ clknet_leaf_12_CLK _03786_ VGND VGND VPWR VPWR registers\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32884_ clknet_leaf_351_CLK _00998_ VGND VGND VPWR VPWR registers\[54\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34623_ clknet_leaf_189_CLK _02737_ VGND VGND VPWR VPWR registers\[27\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31835_ _09676_ registers\[49\]\[9\] _14419_ VGND VGND VPWR VPWR _14429_ sky130_fd_sc_hd__mux2_1
X_19557_ registers\[16\]\[33\] registers\[17\]\[33\] registers\[18\]\[33\] registers\[19\]\[33\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__mux4_1
X_16769_ _14991_ _15261_ _15262_ _14996_ VGND VGND VPWR VPWR _15263_ sky130_fd_sc_hd__a22o_1
XFILLER_111_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18508_ _05197_ _05265_ _05266_ _05202_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__a22o_1
XFILLER_55_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34554_ clknet_leaf_184_CLK _02668_ VGND VGND VPWR VPWR registers\[28\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31766_ registers\[59\]\[40\] net35 _14392_ VGND VGND VPWR VPWR _14393_ sky130_fd_sc_hd__mux2_1
XFILLER_202_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19488_ _06182_ _06218_ _06219_ _06185_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__a22o_1
XFILLER_34_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30717_ registers\[12\]\[55\] _13050_ _13835_ VGND VGND VPWR VPWR _13841_ sky130_fd_sc_hd__mux2_1
XFILLER_210_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33505_ clknet_leaf_35_CLK _01619_ VGND VGND VPWR VPWR registers\[44\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_18439_ registers\[40\]\[2\] registers\[41\]\[2\] registers\[42\]\[2\] registers\[43\]\[2\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31697_ _14356_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__clkbuf_1
X_34485_ clknet_leaf_414_CLK _02599_ VGND VGND VPWR VPWR registers\[2\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36224_ clknet_leaf_117_CLK _00109_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dfxtp_1
X_21450_ registers\[44\]\[22\] registers\[45\]\[22\] registers\[46\]\[22\] registers\[47\]\[22\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__mux4_1
X_33436_ clknet_leaf_30_CLK _01550_ VGND VGND VPWR VPWR registers\[45\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_30648_ registers\[12\]\[22\] _12981_ _13802_ VGND VGND VPWR VPWR _13805_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20401_ _07102_ _07105_ _06847_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__o21ba_2
XFILLER_120_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33367_ clknet_leaf_123_CLK _01481_ VGND VGND VPWR VPWR registers\[46\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_36155_ clknet_leaf_282_CLK _04269_ VGND VGND VPWR VPWR registers\[49\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21381_ registers\[52\]\[20\] registers\[53\]\[20\] registers\[54\]\[20\] registers\[55\]\[20\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__mux4_1
X_30579_ _13768_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20332_ _07036_ _07039_ _06880_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__o21ba_1
X_23120_ _09680_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
X_35106_ clknet_leaf_466_CLK _03220_ VGND VGND VPWR VPWR registers\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_32318_ clknet_leaf_191_CLK _00432_ VGND VGND VPWR VPWR registers\[19\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_33298_ clknet_leaf_123_CLK _01412_ VGND VGND VPWR VPWR registers\[47\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_36086_ clknet_leaf_328_CLK _04200_ VGND VGND VPWR VPWR registers\[59\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23051_ _09630_ registers\[62\]\[55\] _09620_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__mux2_1
X_20263_ registers\[16\]\[53\] registers\[17\]\[53\] registers\[18\]\[53\] registers\[19\]\[53\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__mux4_1
X_32249_ clknet_leaf_281_CLK _00363_ VGND VGND VPWR VPWR registers\[39\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_35037_ clknet_leaf_491_CLK _03151_ VGND VGND VPWR VPWR registers\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22002_ registers\[32\]\[38\] registers\[33\]\[38\] registers\[34\]\[38\] registers\[35\]\[38\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__mux4_1
XTAP_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20194_ _06868_ _06904_ _06905_ _06871_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__a22o_1
XFILLER_62_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26810_ _11722_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__clkbuf_1
XTAP_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27790_ registers\[33\]\[43\] _10395_ _12266_ VGND VGND VPWR VPWR _12270_ sky130_fd_sc_hd__mux2_1
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26741_ _11686_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23953_ _10149_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35939_ clknet_leaf_470_CLK _04053_ VGND VGND VPWR VPWR registers\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22904_ net63 VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__clkbuf_4
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29460_ _13179_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__clkbuf_1
X_26672_ _11649_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__clkbuf_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23884_ _10113_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_905 _09662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28411_ _12596_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_1
X_25623_ _11096_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_916 _09756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22835_ _09468_ _09471_ _07369_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__o21ba_1
X_29391_ _13143_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_927 _09869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_938 _10232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_949 _10410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28342_ registers\[2\]\[49\] _10407_ _12550_ VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__mux2_1
X_25554_ registers\[4\]\[42\] _10393_ _11056_ VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__mux2_1
XFILLER_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22766_ registers\[52\]\[60\] registers\[53\]\[60\] registers\[54\]\[60\] registers\[55\]\[60\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__mux4_1
XFILLER_112_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ _10471_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28273_ registers\[2\]\[16\] _10338_ _12517_ VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__mux2_1
X_21717_ _08383_ _08386_ _08087_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__o21ba_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25485_ _11022_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22697_ _09148_ _09336_ _09337_ _09153_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__a22o_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27224_ _11971_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__clkbuf_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24436_ _10433_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
X_21648_ registers\[40\]\[28\] registers\[41\]\[28\] registers\[42\]\[28\] registers\[43\]\[28\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__mux4_1
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27155_ _11934_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_193_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_193_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24367_ registers\[57\]\[39\] _10386_ _10368_ VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21579_ registers\[32\]\[26\] registers\[33\]\[26\] registers\[34\]\[26\] registers\[35\]\[26\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__mux4_1
XANTENNA_91 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26106_ _11351_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
X_23318_ _09807_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27086_ _11792_ registers\[38\]\[30\] _11898_ VGND VGND VPWR VPWR _11899_ sky130_fd_sc_hd__mux2_1
X_24298_ net9 VGND VGND VPWR VPWR _10340_ sky130_fd_sc_hd__buf_4
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26037_ _11315_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23249_ _09761_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1304 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1315 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1326 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17810_ registers\[8\]\[49\] registers\[9\]\[49\] registers\[10\]\[49\] registers\[11\]\[49\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__mux4_1
XANTENNA_1337 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1348 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18790_ _05042_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__buf_4
XTAP_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27988_ _11748_ registers\[31\]\[9\] _12364_ VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__mux2_1
XANTENNA_1359 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ registers\[12\]\[47\] registers\[13\]\[47\] registers\[14\]\[47\] registers\[15\]\[47\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux4_1
XFILLER_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29727_ registers\[1\]\[34\] _13006_ _13315_ VGND VGND VPWR VPWR _13320_ sky130_fd_sc_hd__mux2_1
X_26939_ _11808_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_1
XTAP_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17672_ registers\[4\]\[45\] registers\[5\]\[45\] registers\[6\]\[45\] registers\[7\]\[45\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__mux4_1
X_29658_ registers\[1\]\[1\] _12937_ _13282_ VGND VGND VPWR VPWR _13284_ sky130_fd_sc_hd__mux2_1
XFILLER_78_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16623_ _15098_ _15105_ _15114_ _15121_ VGND VGND VPWR VPWR _15122_ sky130_fd_sc_hd__or4_1
X_19411_ registers\[24\]\[29\] registers\[25\]\[29\] registers\[26\]\[29\] registers\[27\]\[29\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__mux4_1
XFILLER_210_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28609_ _12700_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29589_ _13247_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31620_ registers\[63\]\[35\] net29 _14310_ VGND VGND VPWR VPWR _14316_ sky130_fd_sc_hd__mux2_1
X_16554_ registers\[20\]\[13\] registers\[21\]\[13\] registers\[22\]\[13\] registers\[23\]\[13\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15055_ sky130_fd_sc_hd__mux4_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19342_ registers\[28\]\[27\] registers\[29\]\[27\] registers\[30\]\[27\] registers\[31\]\[27\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__mux4_1
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31551_ registers\[63\]\[2\] net23 _14277_ VGND VGND VPWR VPWR _14280_ sky130_fd_sc_hd__mux2_1
X_19273_ registers\[20\]\[25\] registers\[21\]\[25\] registers\[22\]\[25\] registers\[23\]\[25\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16485_ _14952_ _14986_ _14987_ _14957_ VGND VGND VPWR VPWR _14988_ sky130_fd_sc_hd__a22o_1
XFILLER_188_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18224_ _14587_ _04987_ _04988_ _14597_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a22o_1
X_30502_ _09693_ registers\[13\]\[17\] _13720_ VGND VGND VPWR VPWR _13728_ sky130_fd_sc_hd__mux2_1
XFILLER_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34270_ clknet_leaf_22_CLK _02384_ VGND VGND VPWR VPWR registers\[32\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31482_ _14243_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33221_ clknet_leaf_232_CLK _01335_ VGND VGND VPWR VPWR registers\[4\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18155_ registers\[40\]\[60\] registers\[41\]\[60\] registers\[42\]\[60\] registers\[43\]\[60\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__mux4_1
X_30433_ _13691_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_184_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_184_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17106_ _15482_ _15589_ _15590_ _15485_ VGND VGND VPWR VPWR _15591_ sky130_fd_sc_hd__a22o_1
X_33152_ clknet_leaf_269_CLK _01266_ VGND VGND VPWR VPWR registers\[50\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18086_ registers\[24\]\[57\] registers\[25\]\[57\] registers\[26\]\[57\] registers\[27\]\[57\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__mux4_1
XFILLER_172_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30364_ _13655_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32103_ clknet_leaf_483_CLK _00017_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17037_ _15487_ _15522_ _15523_ _15490_ VGND VGND VPWR VPWR _15524_ sky130_fd_sc_hd__a22o_1
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33083_ clknet_leaf_285_CLK _01197_ VGND VGND VPWR VPWR registers\[51\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_30295_ _13618_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__clkbuf_1
X_32034_ clknet_leaf_445_CLK _00212_ VGND VGND VPWR VPWR registers\[62\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18988_ _05496_ _05732_ _05733_ _05499_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__a22o_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17939_ registers\[40\]\[53\] registers\[41\]\[53\] registers\[42\]\[53\] registers\[43\]\[53\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux4_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33985_ clknet_leaf_258_CLK _02099_ VGND VGND VPWR VPWR registers\[37\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35724_ clknet_leaf_144_CLK _03838_ VGND VGND VPWR VPWR registers\[10\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_20950_ _07316_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__buf_4
X_32936_ clknet_leaf_423_CLK _01050_ VGND VGND VPWR VPWR registers\[53\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19609_ registers\[60\]\[35\] registers\[61\]\[35\] registers\[62\]\[35\] registers\[63\]\[35\]
+ _06305_ _06099_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__mux4_1
XFILLER_26_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35655_ clknet_leaf_216_CLK _03769_ VGND VGND VPWR VPWR registers\[11\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20881_ _07313_ _07572_ _07573_ _07322_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__a22o_1
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32867_ clknet_leaf_443_CLK _00981_ VGND VGND VPWR VPWR registers\[54\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22620_ registers\[0\]\[55\] registers\[1\]\[55\] registers\[2\]\[55\] registers\[3\]\[55\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__mux4_1
X_34606_ clknet_leaf_410_CLK _02720_ VGND VGND VPWR VPWR registers\[27\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_31818_ _14420_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35586_ clknet_leaf_238_CLK _03700_ VGND VGND VPWR VPWR registers\[12\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32798_ clknet_leaf_46_CLK _00912_ VGND VGND VPWR VPWR registers\[55\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22551_ _09020_ _09195_ _09196_ _09024_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__a22o_1
X_34537_ clknet_leaf_404_CLK _02651_ VGND VGND VPWR VPWR registers\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31749_ registers\[59\]\[32\] net26 _14381_ VGND VGND VPWR VPWR _14384_ sky130_fd_sc_hd__mux2_1
XFILLER_195_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21502_ _08172_ _08177_ _08073_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25270_ _10810_ registers\[51\]\[38\] _10898_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__mux2_1
X_22482_ registers\[52\]\[51\] registers\[53\]\[51\] registers\[54\]\[51\] registers\[55\]\[51\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__mux4_1
X_34468_ clknet_leaf_464_CLK _02582_ VGND VGND VPWR VPWR registers\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24221_ _10291_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
X_36207_ clknet_leaf_100_CLK _00090_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dfxtp_1
X_33419_ clknet_leaf_164_CLK _01533_ VGND VGND VPWR VPWR registers\[46\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21433_ registers\[24\]\[21\] registers\[25\]\[21\] registers\[26\]\[21\] registers\[27\]\[21\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_175_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_175_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34399_ clknet_leaf_488_CLK _02513_ VGND VGND VPWR VPWR registers\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21364_ _08040_ _08043_ _07744_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24152_ _10232_ VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__buf_4
X_36138_ clknet_leaf_425_CLK _04252_ VGND VGND VPWR VPWR registers\[49\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23103_ registers\[39\]\[5\] _09668_ _09658_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__mux2_1
X_20315_ registers\[60\]\[55\] registers\[61\]\[55\] registers\[62\]\[55\] registers\[63\]\[55\]
+ _06991_ _06785_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__mux4_1
XFILLER_159_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24083_ _10218_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28960_ _12885_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__clkbuf_1
X_36069_ clknet_leaf_438_CLK _04183_ VGND VGND VPWR VPWR registers\[59\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_21295_ registers\[40\]\[18\] registers\[41\]\[18\] registers\[42\]\[18\] registers\[43\]\[18\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__mux4_1
XFILLER_239_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23034_ net46 VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__buf_4
X_20246_ registers\[56\]\[53\] registers\[57\]\[53\] registers\[58\]\[53\] registers\[59\]\[53\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__mux4_1
X_27911_ _12333_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__clkbuf_1
X_28891_ _11841_ registers\[25\]\[53\] _12845_ VGND VGND VPWR VPWR _12849_ sky130_fd_sc_hd__mux2_1
XFILLER_235_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27842_ _12297_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__clkbuf_1
X_20177_ _06885_ _06888_ _06847_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__o21ba_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27773_ registers\[33\]\[35\] _10378_ _12255_ VGND VGND VPWR VPWR _12261_ sky130_fd_sc_hd__mux2_1
X_24985_ _09644_ registers\[53\]\[62\] _10657_ VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__mux2_1
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29512_ _13206_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__clkbuf_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26724_ _11677_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _10140_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_702 _07278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29443_ _13170_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26655_ _11640_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_713 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23867_ _10104_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_724 _07344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_735 _07356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_746 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25606_ registers\[48\]\[1\] _10307_ _11086_ VGND VGND VPWR VPWR _11088_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29374_ _09817_ registers\[22\]\[59\] _13124_ VGND VGND VPWR VPWR _13134_ sky130_fd_sc_hd__mux2_1
XFILLER_199_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22818_ registers\[44\]\[62\] registers\[45\]\[62\] registers\[46\]\[62\] registers\[47\]\[62\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__mux4_1
XANTENNA_757 _07388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26586_ _11604_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_1
X_23798_ _10067_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_768 _07687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_779 _08318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28325_ _12551_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25537_ registers\[4\]\[34\] _10376_ _11045_ VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__mux2_1
X_22749_ registers\[28\]\[59\] registers\[29\]\[59\] registers\[30\]\[59\] registers\[31\]\[59\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__mux4_1
XFILLER_158_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16270_ _14755_ _14762_ _14771_ _14778_ VGND VGND VPWR VPWR _14779_ sky130_fd_sc_hd__or4_2
X_28256_ registers\[2\]\[8\] _10321_ _12506_ VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__mux2_1
X_25468_ registers\[4\]\[1\] _10307_ _11012_ VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_52__f_CLK clknet_5_26_0_CLK VGND VGND VPWR VPWR clknet_6_52__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_27207_ _11962_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__clkbuf_1
X_24419_ net52 VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__buf_4
XFILLER_200_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_166_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_166_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28187_ _12478_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25399_ _10975_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__clkbuf_1
X_27138_ _11845_ registers\[38\]\[55\] _11920_ VGND VGND VPWR VPWR _11926_ sky130_fd_sc_hd__mux2_1
XFILLER_181_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19960_ registers\[48\]\[45\] registers\[49\]\[45\] registers\[50\]\[45\] registers\[51\]\[45\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__mux4_1
X_27069_ _11776_ registers\[38\]\[22\] _11887_ VGND VGND VPWR VPWR _11890_ sky130_fd_sc_hd__mux2_1
XFILLER_181_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18911_ _05345_ _05657_ _05658_ _05348_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a22o_1
XFILLER_84_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30080_ _13505_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__clkbuf_1
XTAP_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19891_ _06576_ _06609_ _06610_ _06579_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__a22o_1
XTAP_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1101 _14530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1112 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1123 _14578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18842_ registers\[0\]\[13\] registers\[1\]\[13\] registers\[2\]\[13\] registers\[3\]\[13\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__mux4_1
XFILLER_45_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1134 _14610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1145 _15245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1156 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1167 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1178 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15985_ net67 net68 VGND VGND VPWR VPWR _14499_ sky130_fd_sc_hd__nor2_4
X_18773_ registers\[8\]\[11\] registers\[9\]\[11\] registers\[10\]\[11\] registers\[11\]\[11\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__mux4_1
XFILLER_62_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1189 _15845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17724_ _04333_ _04502_ _04503_ _04338_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__a22o_1
XFILLER_23_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30982_ _13980_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33770_ clknet_leaf_427_CLK _01884_ VGND VGND VPWR VPWR registers\[40\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32721_ clknet_leaf_72_CLK _00835_ VGND VGND VPWR VPWR registers\[56\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17655_ registers\[44\]\[45\] registers\[45\]\[45\] registers\[46\]\[45\] registers\[47\]\[45\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux4_1
XFILLER_35_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35440_ clknet_leaf_375_CLK _03554_ VGND VGND VPWR VPWR registers\[14\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16606_ _15101_ _15104_ _14934_ _14935_ VGND VGND VPWR VPWR _15105_ sky130_fd_sc_hd__o211a_2
X_32652_ clknet_leaf_167_CLK _00766_ VGND VGND VPWR VPWR registers\[58\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_17586_ registers\[40\]\[43\] registers\[41\]\[43\] registers\[42\]\[43\] registers\[43\]\[43\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__mux4_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16537_ registers\[60\]\[13\] registers\[61\]\[13\] registers\[62\]\[13\] registers\[63\]\[13\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _15038_ sky130_fd_sc_hd__mux4_1
X_31603_ registers\[63\]\[27\] net20 _14299_ VGND VGND VPWR VPWR _14307_ sky130_fd_sc_hd__mux2_1
X_19325_ registers\[56\]\[27\] registers\[57\]\[27\] registers\[58\]\[27\] registers\[59\]\[27\]
+ _05958_ _05748_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__mux4_1
X_32583_ clknet_leaf_210_CLK _00697_ VGND VGND VPWR VPWR registers\[5\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35371_ clknet_leaf_397_CLK _03485_ VGND VGND VPWR VPWR registers\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34322_ clknet_leaf_99_CLK _02436_ VGND VGND VPWR VPWR registers\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_31534_ _14270_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16468_ _14855_ _14969_ _14970_ _14861_ VGND VGND VPWR VPWR _14971_ sky130_fd_sc_hd__a22o_1
X_19256_ registers\[60\]\[25\] registers\[61\]\[25\] registers\[62\]\[25\] registers\[63\]\[25\]
+ _05962_ _05756_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__mux4_1
XFILLER_143_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18207_ registers\[16\]\[61\] registers\[17\]\[61\] registers\[18\]\[61\] registers\[19\]\[61\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__mux4_1
XFILLER_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_157_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_157_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34253_ clknet_leaf_76_CLK _02367_ VGND VGND VPWR VPWR registers\[33\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_31465_ _14234_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__clkbuf_1
X_19187_ registers\[56\]\[23\] registers\[57\]\[23\] registers\[58\]\[23\] registers\[59\]\[23\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__mux4_1
X_16399_ registers\[0\]\[9\] registers\[1\]\[9\] registers\[2\]\[9\] registers\[3\]\[9\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14904_ sky130_fd_sc_hd__mux4_1
X_18138_ _04902_ _04905_ _04619_ _04620_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__o211a_1
X_33204_ clknet_leaf_321_CLK _01318_ VGND VGND VPWR VPWR registers\[4\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30416_ _09775_ registers\[14\]\[40\] _13682_ VGND VGND VPWR VPWR _13683_ sky130_fd_sc_hd__mux2_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34184_ clknet_leaf_244_CLK _02298_ VGND VGND VPWR VPWR registers\[34\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31396_ registers\[7\]\[57\] net53 _14190_ VGND VGND VPWR VPWR _14198_ sky130_fd_sc_hd__mux2_1
XFILLER_144_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18069_ registers\[36\]\[57\] registers\[37\]\[57\] registers\[38\]\[57\] registers\[39\]\[57\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30347_ _13646_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__clkbuf_1
X_33135_ clknet_leaf_365_CLK _01249_ VGND VGND VPWR VPWR registers\[50\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20100_ registers\[36\]\[49\] registers\[37\]\[49\] registers\[38\]\[49\] registers\[39\]\[49\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1078 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21080_ registers\[24\]\[11\] registers\[25\]\[11\] registers\[26\]\[11\] registers\[27\]\[11\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__mux4_1
X_33066_ clknet_leaf_419_CLK _01180_ VGND VGND VPWR VPWR registers\[51\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_30278_ _13609_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32017_ clknet_leaf_179_CLK _00195_ VGND VGND VPWR VPWR registers\[62\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_20031_ registers\[56\]\[47\] registers\[57\]\[47\] registers\[58\]\[47\] registers\[59\]\[47\]
+ _06644_ _06434_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__mux4_1
XFILLER_8_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1690 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24770_ _10613_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33968_ clknet_leaf_357_CLK _02082_ VGND VGND VPWR VPWR registers\[37\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_21982_ registers\[52\]\[37\] registers\[53\]\[37\] registers\[54\]\[37\] registers\[55\]\[37\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__mux4_1
XFILLER_230_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _09533_ registers\[29\]\[9\] _10017_ VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__mux2_1
X_35707_ clknet_leaf_301_CLK _03821_ VGND VGND VPWR VPWR registers\[10\]\[45\] sky130_fd_sc_hd__dfxtp_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20933_ registers\[24\]\[7\] registers\[25\]\[7\] registers\[26\]\[7\] registers\[27\]\[7\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__mux4_1
X_32919_ clknet_leaf_63_CLK _01033_ VGND VGND VPWR VPWR registers\[53\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33899_ clknet_leaf_424_CLK _02013_ VGND VGND VPWR VPWR registers\[38\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26440_ _11527_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__clkbuf_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35638_ clknet_leaf_330_CLK _03752_ VGND VGND VPWR VPWR registers\[11\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_23652_ _09989_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
X_20864_ registers\[16\]\[5\] registers\[17\]\[5\] registers\[18\]\[5\] registers\[19\]\[5\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__mux4_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22603_ _09222_ _09231_ _09238_ _09247_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__or4_4
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26371_ _10821_ registers\[43\]\[43\] _11487_ VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__mux2_1
X_23583_ registers\[61\]\[9\] _09676_ _09943_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_396_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_396_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35569_ clknet_leaf_380_CLK _03683_ VGND VGND VPWR VPWR registers\[12\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20795_ _07355_ _07489_ _07490_ _07367_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__a22o_1
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28110_ _12438_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25322_ _10862_ registers\[51\]\[63\] _10864_ VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__mux2_1
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22534_ registers\[20\]\[52\] registers\[21\]\[52\] registers\[22\]\[52\] registers\[23\]\[52\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__mux4_1
X_29090_ registers\[23\]\[12\] _12960_ _12956_ VGND VGND VPWR VPWR _12961_ sky130_fd_sc_hd__mux2_1
XFILLER_183_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28041_ _11801_ registers\[31\]\[34\] _12397_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25253_ _10864_ VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_148_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_148_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22465_ _07366_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24204_ _10282_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_21416_ registers\[36\]\[21\] registers\[37\]\[21\] registers\[38\]\[21\] registers\[39\]\[21\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__mux4_1
X_25184_ _10860_ registers\[52\]\[62\] _10730_ VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__mux2_1
X_22396_ _07289_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__buf_4
X_24135_ _10246_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21347_ registers\[60\]\[19\] registers\[61\]\[19\] registers\[62\]\[19\] registers\[63\]\[19\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__mux4_1
X_29992_ _13459_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24066_ _10209_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__clkbuf_1
X_28943_ _12876_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21278_ _07956_ _07959_ _07719_ _07720_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__o211a_1
X_23017_ _09607_ registers\[62\]\[44\] _09599_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__mux2_1
X_20229_ registers\[16\]\[52\] registers\[17\]\[52\] registers\[18\]\[52\] registers\[19\]\[52\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_320_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_320_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28874_ _11824_ registers\[25\]\[45\] _12834_ VGND VGND VPWR VPWR _12840_ sky130_fd_sc_hd__mux2_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27825_ registers\[33\]\[60\] _10430_ _12221_ VGND VGND VPWR VPWR _12288_ sky130_fd_sc_hd__mux2_1
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24968_ _10717_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27756_ registers\[33\]\[27\] _10361_ _12244_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__mux2_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26707_ _11668_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23919_ _10131_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
X_27687_ _12215_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__clkbuf_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24899_ _10681_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_510 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_217_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_521 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_532 _00176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _15915_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__clkbuf_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29426_ _13161_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26638_ _10817_ registers\[41\]\[41\] _11630_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__mux2_1
XANTENNA_543 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_554 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_565 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_576 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _15677_ _15846_ _15847_ _15682_ VGND VGND VPWR VPWR _15848_ sky130_fd_sc_hd__a22o_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_587 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26569_ _11595_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__clkbuf_1
X_29357_ _13125_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_387_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_387_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_598 _05088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16322_ registers\[60\]\[7\] registers\[61\]\[7\] registers\[62\]\[7\] registers\[63\]\[7\]
+ _14727_ _14544_ VGND VGND VPWR VPWR _14829_ sky130_fd_sc_hd__mux4_1
X_19110_ _05819_ _05828_ _05838_ _05852_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__or4_4
XFILLER_213_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28308_ _12542_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__clkbuf_1
X_29288_ _09695_ registers\[22\]\[18\] _13080_ VGND VGND VPWR VPWR _13089_ sky130_fd_sc_hd__mux2_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19041_ registers\[36\]\[19\] registers\[37\]\[19\] registers\[38\]\[19\] registers\[39\]\[19\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__mux4_1
X_28239_ _12505_ VGND VGND VPWR VPWR _12506_ sky130_fd_sc_hd__buf_4
X_16253_ _14758_ _14761_ _14554_ _14556_ VGND VGND VPWR VPWR _14762_ sky130_fd_sc_hd__o211a_1
XFILLER_146_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_139_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_139_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31250_ _14121_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__clkbuf_1
X_16184_ registers\[60\]\[3\] registers\[61\]\[3\] registers\[62\]\[3\] registers\[63\]\[3\]
+ _14542_ _14544_ VGND VGND VPWR VPWR _14695_ sky130_fd_sc_hd__mux4_1
XFILLER_51_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30201_ _13569_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput208 net208 VGND VGND VPWR VPWR D2[59] sky130_fd_sc_hd__buf_2
XFILLER_177_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31181_ registers\[8\]\[19\] net11 _14075_ VGND VGND VPWR VPWR _14085_ sky130_fd_sc_hd__mux2_1
Xoutput219 net219 VGND VGND VPWR VPWR D3[10] sky130_fd_sc_hd__buf_2
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30132_ registers\[16\]\[34\] _13006_ _13528_ VGND VGND VPWR VPWR _13533_ sky130_fd_sc_hd__mux2_1
X_19943_ registers\[24\]\[44\] registers\[25\]\[44\] registers\[26\]\[44\] registers\[27\]\[44\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux4_1
XFILLER_142_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30063_ registers\[16\]\[1\] _12937_ _13495_ VGND VGND VPWR VPWR _13497_ sky130_fd_sc_hd__mux2_1
X_34940_ clknet_leaf_307_CLK _03054_ VGND VGND VPWR VPWR registers\[22\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_19874_ _06591_ _06594_ _06523_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_311_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_311_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18825_ _05552_ _05559_ _05566_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__or4_2
XTAP_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34871_ clknet_leaf_308_CLK _02985_ VGND VGND VPWR VPWR registers\[23\]\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33822_ clknet_leaf_487_CLK _01936_ VGND VGND VPWR VPWR registers\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18756_ _05500_ _05507_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__o21ba_1
XFILLER_237_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17707_ registers\[4\]\[46\] registers\[5\]\[46\] registers\[6\]\[46\] registers\[7\]\[46\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__mux4_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33753_ clknet_leaf_90_CLK _01867_ VGND VGND VPWR VPWR registers\[40\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18687_ registers\[44\]\[9\] registers\[45\]\[9\] registers\[46\]\[9\] registers\[47\]\[9\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__mux4_1
X_30965_ _13971_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32704_ clknet_leaf_267_CLK _00818_ VGND VGND VPWR VPWR registers\[57\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_17638_ registers\[4\]\[44\] registers\[5\]\[44\] registers\[6\]\[44\] registers\[7\]\[44\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__mux4_1
XFILLER_97_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33684_ clknet_leaf_119_CLK _01798_ VGND VGND VPWR VPWR registers\[41\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30896_ _13935_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__clkbuf_1
X_35423_ clknet_leaf_482_CLK _03537_ VGND VGND VPWR VPWR registers\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32635_ clknet_leaf_284_CLK _00749_ VGND VGND VPWR VPWR registers\[58\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_17569_ registers\[0\]\[42\] registers\[1\]\[42\] registers\[2\]\[42\] registers\[3\]\[42\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_378_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_378_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19308_ registers\[16\]\[26\] registers\[17\]\[26\] registers\[18\]\[26\] registers\[19\]\[26\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__mux4_1
XFILLER_225_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20580_ _07278_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__buf_6
XFILLER_17_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35354_ clknet_leaf_13_CLK _03468_ VGND VGND VPWR VPWR registers\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32566_ clknet_leaf_319_CLK _00680_ VGND VGND VPWR VPWR registers\[5\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34305_ clknet_leaf_257_CLK _02419_ VGND VGND VPWR VPWR registers\[32\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31517_ _09797_ registers\[6\]\[50\] _14261_ VGND VGND VPWR VPWR _14262_ sky130_fd_sc_hd__mux2_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19239_ _05839_ _05976_ _05977_ _05842_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__a22o_1
XFILLER_165_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35285_ clknet_leaf_89_CLK _03399_ VGND VGND VPWR VPWR registers\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32497_ clknet_leaf_367_CLK _00611_ VGND VGND VPWR VPWR registers\[60\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_34236_ clknet_leaf_276_CLK _02350_ VGND VGND VPWR VPWR registers\[33\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_22250_ _08879_ _08888_ _08895_ _08904_ VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__or4_4
XFILLER_180_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31448_ _14225_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21201_ registers\[48\]\[15\] registers\[49\]\[15\] registers\[50\]\[15\] registers\[51\]\[15\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22181_ registers\[20\]\[42\] registers\[21\]\[42\] registers\[22\]\[42\] registers\[23\]\[42\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__mux4_1
X_31379_ registers\[7\]\[49\] net44 _14179_ VGND VGND VPWR VPWR _14189_ sky130_fd_sc_hd__mux2_1
X_34167_ clknet_leaf_342_CLK _02281_ VGND VGND VPWR VPWR registers\[34\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21132_ _07783_ _07816_ _07817_ _07786_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__a22o_1
X_33118_ clknet_leaf_37_CLK _01232_ VGND VGND VPWR VPWR registers\[50\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_34098_ clknet_leaf_355_CLK _02212_ VGND VGND VPWR VPWR registers\[35\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21063_ registers\[36\]\[11\] registers\[37\]\[11\] registers\[38\]\[11\] registers\[39\]\[11\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__mux4_1
X_25940_ _11264_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_302_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_302_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33049_ clknet_leaf_35_CLK _01163_ VGND VGND VPWR VPWR registers\[51\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20014_ registers\[16\]\[46\] registers\[17\]\[46\] registers\[18\]\[46\] registers\[19\]\[46\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__mux4_1
XFILLER_63_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25871_ _11227_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24822_ _10640_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27610_ _12175_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28590_ _12690_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__clkbuf_1
X_27541_ _11843_ registers\[35\]\[54\] _12133_ VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24753_ _10604_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__clkbuf_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _08423_ _08626_ _08627_ _08428_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__a22o_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _10018_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ registers\[36\]\[7\] registers\[37\]\[7\] registers\[38\]\[7\] registers\[39\]\[7\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__mux4_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27472_ _11774_ registers\[35\]\[21\] _12100_ VGND VGND VPWR VPWR _12102_ sky130_fd_sc_hd__mux2_1
X_24684_ _09615_ registers\[55\]\[48\] _10558_ VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__mux2_1
XFILLER_203_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21896_ _08557_ _08560_ _08430_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__o21ba_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26423_ _11518_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29211_ registers\[23\]\[51\] _13042_ _13040_ VGND VGND VPWR VPWR _13043_ sky130_fd_sc_hd__mux2_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23635_ _09980_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ registers\[56\]\[5\] registers\[57\]\[5\] registers\[58\]\[5\] registers\[59\]\[5\]
+ _07508_ _07317_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__mux4_1
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_369_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_369_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29142_ registers\[23\]\[29\] _12995_ _12977_ VGND VGND VPWR VPWR _12996_ sky130_fd_sc_hd__mux2_1
X_26354_ _10804_ registers\[43\]\[35\] _11476_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__mux2_1
X_23566_ _09944_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
X_20778_ registers\[36\]\[3\] registers\[37\]\[3\] registers\[38\]\[3\] registers\[39\]\[3\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__mux4_1
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25305_ _10925_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22517_ registers\[60\]\[52\] registers\[61\]\[52\] registers\[62\]\[52\] registers\[63\]\[52\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__mux4_1
X_29073_ net62 VGND VGND VPWR VPWR _12949_ sky130_fd_sc_hd__clkbuf_4
X_26285_ _10735_ registers\[43\]\[2\] _11443_ VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__mux2_1
X_23497_ _09584_ registers\[19\]\[33\] _09903_ VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__mux2_1
X_28024_ _11784_ registers\[31\]\[26\] _12386_ VGND VGND VPWR VPWR _12393_ sky130_fd_sc_hd__mux2_1
XFILLER_167_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25236_ _10889_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__clkbuf_1
X_22448_ registers\[0\]\[50\] registers\[1\]\[50\] registers\[2\]\[50\] registers\[3\]\[50\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__mux4_1
XFILLER_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25167_ _10849_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22379_ registers\[12\]\[48\] registers\[13\]\[48\] registers\[14\]\[48\] registers\[15\]\[48\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__mux4_1
XFILLER_108_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24118_ _10237_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25098_ _10802_ registers\[52\]\[34\] _10794_ VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__mux2_1
X_29975_ _13450_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28926_ _12867_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24049_ _10200_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__clkbuf_1
X_16940_ registers\[28\]\[24\] registers\[29\]\[24\] registers\[30\]\[24\] registers\[31\]\[24\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15430_ sky130_fd_sc_hd__mux4_1
XFILLER_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16871_ _15290_ _15361_ _15362_ _15293_ VGND VGND VPWR VPWR _15363_ sky130_fd_sc_hd__a22o_1
X_28857_ _11807_ registers\[25\]\[37\] _12823_ VGND VGND VPWR VPWR _12831_ sky130_fd_sc_hd__mux2_1
X_18610_ registers\[40\]\[7\] registers\[41\]\[7\] registers\[42\]\[7\] registers\[43\]\[7\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__mux4_1
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27808_ _12279_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__clkbuf_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ registers\[24\]\[34\] registers\[25\]\[34\] registers\[26\]\[34\] registers\[27\]\[34\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__mux4_1
XFILLER_219_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28788_ _11738_ registers\[25\]\[4\] _12790_ VGND VGND VPWR VPWR _12795_ sky130_fd_sc_hd__mux2_1
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18541_ registers\[32\]\[5\] registers\[33\]\[5\] registers\[34\]\[5\] registers\[35\]\[5\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__mux4_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27739_ registers\[33\]\[19\] _10344_ _12233_ VGND VGND VPWR VPWR _12243_ sky130_fd_sc_hd__mux2_1
XFILLER_92_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _05209_ _05216_ _05223_ _05232_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__or4_4
X_30750_ _13858_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29409_ _09681_ registers\[21\]\[11\] _13151_ VGND VGND VPWR VPWR _13153_ sky130_fd_sc_hd__mux2_1
X_17423_ registers\[8\]\[38\] registers\[9\]\[38\] registers\[10\]\[38\] registers\[11\]\[38\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15899_ sky130_fd_sc_hd__mux4_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_373 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30681_ registers\[12\]\[38\] _13014_ _13813_ VGND VGND VPWR VPWR _13822_ sky130_fd_sc_hd__mux2_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32420_ clknet_leaf_472_CLK _00534_ VGND VGND VPWR VPWR registers\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17354_ registers\[4\]\[36\] registers\[5\]\[36\] registers\[6\]\[36\] registers\[7\]\[36\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15832_ sky130_fd_sc_hd__mux4_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16305_ registers\[20\]\[6\] registers\[21\]\[6\] registers\[22\]\[6\] registers\[23\]\[6\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14813_ sky130_fd_sc_hd__mux4_1
XFILLER_146_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17285_ registers\[4\]\[34\] registers\[5\]\[34\] registers\[6\]\[34\] registers\[7\]\[34\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15765_ sky130_fd_sc_hd__mux4_1
X_32351_ clknet_leaf_50_CLK _00465_ VGND VGND VPWR VPWR registers\[61\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16236_ _14601_ _14744_ _14745_ _14611_ VGND VGND VPWR VPWR _14746_ sky130_fd_sc_hd__a22o_1
X_19024_ _05693_ _05765_ _05768_ _05696_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__a22o_1
X_31302_ registers\[7\]\[12\] net4 _14146_ VGND VGND VPWR VPWR _14149_ sky130_fd_sc_hd__mux2_1
X_35070_ clknet_leaf_188_CLK _03184_ VGND VGND VPWR VPWR registers\[20\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_32282_ clknet_leaf_20_CLK _00396_ VGND VGND VPWR VPWR registers\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31233_ _14112_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__clkbuf_1
X_34021_ clknet_leaf_433_CLK _02135_ VGND VGND VPWR VPWR registers\[36\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_983 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16167_ _14603_ VGND VGND VPWR VPWR _14679_ sky130_fd_sc_hd__buf_6
XFILLER_86_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31164_ _14076_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__clkbuf_1
X_16098_ _14601_ _14605_ _14609_ _14611_ VGND VGND VPWR VPWR _14612_ sky130_fd_sc_hd__a22o_1
XFILLER_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30115_ registers\[16\]\[26\] _12989_ _13517_ VGND VGND VPWR VPWR _13524_ sky130_fd_sc_hd__mux2_1
X_19926_ registers\[56\]\[44\] registers\[57\]\[44\] registers\[58\]\[44\] registers\[59\]\[44\]
+ _06644_ _06434_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__mux4_1
XFILLER_29_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35972_ clknet_leaf_231_CLK _04086_ VGND VGND VPWR VPWR registers\[6\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_31095_ registers\[0\]\[42\] _13023_ _14037_ VGND VGND VPWR VPWR _14040_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30046_ _13487_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34923_ clknet_leaf_458_CLK _03037_ VGND VGND VPWR VPWR registers\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_19857_ registers\[36\]\[42\] registers\[37\]\[42\] registers\[38\]\[42\] registers\[39\]\[42\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__mux4_1
XFILLER_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18808_ _05555_ _05558_ _05483_ _05484_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o211a_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34854_ clknet_leaf_456_CLK _02968_ VGND VGND VPWR VPWR registers\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19788_ _06441_ _06509_ _06510_ _06445_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__a22o_1
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33805_ clknet_leaf_170_CLK _01919_ VGND VGND VPWR VPWR registers\[40\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_18739_ registers\[4\]\[10\] registers\[5\]\[10\] registers\[6\]\[10\] registers\[7\]\[10\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__mux4_1
X_34785_ clknet_leaf_10_CLK _02899_ VGND VGND VPWR VPWR registers\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31997_ clknet_leaf_29_CLK _00169_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33736_ clknet_leaf_243_CLK _01850_ VGND VGND VPWR VPWR registers\[41\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21750_ registers\[24\]\[30\] registers\[25\]\[30\] registers\[26\]\[30\] registers\[27\]\[30\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__mux4_1
X_30948_ _13962_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20701_ _07384_ _07397_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__o21ba_1
X_33667_ clknet_leaf_250_CLK _01781_ VGND VGND VPWR VPWR registers\[42\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21681_ _08075_ _08350_ _08351_ _08078_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__a22o_1
X_30879_ _13926_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__clkbuf_1
X_35406_ clknet_leaf_137_CLK _03520_ VGND VGND VPWR VPWR registers\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_23420_ _09864_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__clkbuf_1
X_20632_ _07277_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__buf_12
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32618_ clknet_leaf_420_CLK _00732_ VGND VGND VPWR VPWR registers\[58\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33598_ clknet_leaf_272_CLK _01712_ VGND VGND VPWR VPWR registers\[43\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35337_ clknet_leaf_155_CLK _03451_ VGND VGND VPWR VPWR registers\[16\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23351_ _09828_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
X_20563_ registers\[4\]\[63\] registers\[5\]\[63\] registers\[6\]\[63\] registers\[7\]\[63\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__mux4_1
X_32549_ clknet_leaf_464_CLK _00663_ VGND VGND VPWR VPWR registers\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22302_ registers\[0\]\[46\] registers\[1\]\[46\] registers\[2\]\[46\] registers\[3\]\[46\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__mux4_1
X_26070_ _11332_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
X_35268_ clknet_leaf_223_CLK _03382_ VGND VGND VPWR VPWR registers\[17\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_23282_ _09783_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20494_ _05136_ _07194_ _07195_ _05146_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__a22o_1
XFILLER_165_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25021_ _10750_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22233_ _08883_ _08887_ _08748_ _08749_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__o211a_1
X_34219_ clknet_leaf_426_CLK _02333_ VGND VGND VPWR VPWR registers\[33\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35199_ clknet_leaf_189_CLK _03313_ VGND VGND VPWR VPWR registers\[18\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22164_ registers\[60\]\[42\] registers\[61\]\[42\] registers\[62\]\[42\] registers\[63\]\[42\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21115_ _07798_ _07801_ _07730_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__o21ba_1
XTAP_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29760_ _13281_ VGND VGND VPWR VPWR _13337_ sky130_fd_sc_hd__buf_4
X_26972_ _11830_ registers\[3\]\[48\] _11814_ VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__mux2_1
X_22095_ registers\[0\]\[40\] registers\[1\]\[40\] registers\[2\]\[40\] registers\[3\]\[40\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__mux4_1
XTAP_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28711_ _12754_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25923_ _11255_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
X_21046_ _07382_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29691_ registers\[1\]\[17\] _12970_ _13293_ VGND VGND VPWR VPWR _13301_ sky130_fd_sc_hd__mux2_1
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28642_ _12717_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__clkbuf_1
X_25854_ _10844_ registers\[47\]\[54\] _11214_ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24805_ _09598_ registers\[54\]\[40\] _10631_ VGND VGND VPWR VPWR _10632_ sky130_fd_sc_hd__mux2_1
X_25785_ _10775_ registers\[47\]\[21\] _11181_ VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__mux2_1
X_28573_ _11792_ registers\[27\]\[30\] _12681_ VGND VGND VPWR VPWR _12682_ sky130_fd_sc_hd__mux2_1
XFILLER_28_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22997_ net32 VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__buf_2
XFILLER_55_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27524_ _11826_ registers\[35\]\[46\] _12122_ VGND VGND VPWR VPWR _12129_ sky130_fd_sc_hd__mux2_1
X_24736_ _10595_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21948_ registers\[8\]\[36\] registers\[9\]\[36\] registers\[10\]\[36\] registers\[11\]\[36\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__mux4_1
XFILLER_83_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27455_ _11757_ registers\[35\]\[13\] _12089_ VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__mux2_1
X_24667_ _10513_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__buf_4
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21879_ _08334_ _08542_ _08543_ _08338_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__a22o_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26406_ _10856_ registers\[43\]\[60\] _11442_ VGND VGND VPWR VPWR _11509_ sky130_fd_sc_hd__mux2_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _09971_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
X_27386_ _12056_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__clkbuf_1
X_24598_ _09529_ registers\[55\]\[7\] _10514_ VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__mux2_1
XFILLER_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26337_ _10787_ registers\[43\]\[27\] _11465_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__mux2_1
X_29125_ _12984_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__clkbuf_1
X_23549_ _09636_ registers\[19\]\[58\] _09925_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__mux2_1
XFILLER_129_939 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29056_ registers\[23\]\[1\] _12937_ _12935_ VGND VGND VPWR VPWR _12938_ sky130_fd_sc_hd__mux2_1
XFILLER_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17070_ registers\[8\]\[28\] registers\[9\]\[28\] registers\[10\]\[28\] registers\[11\]\[28\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15556_ sky130_fd_sc_hd__mux4_1
X_26268_ _11436_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16021_ _14496_ VGND VGND VPWR VPWR _14535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25219_ _10880_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__clkbuf_1
X_28007_ _11767_ registers\[31\]\[18\] _12375_ VGND VGND VPWR VPWR _12384_ sky130_fd_sc_hd__mux2_1
XFILLER_7_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1059 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26199_ _11400_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_70_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_70_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17972_ registers\[32\]\[54\] registers\[33\]\[54\] registers\[34\]\[54\] registers\[35\]\[54\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__mux4_1
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29958_ _13441_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__clkbuf_1
X_19711_ _05090_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__buf_4
X_28909_ _11859_ registers\[25\]\[62\] _12789_ VGND VGND VPWR VPWR _12858_ sky130_fd_sc_hd__mux2_1
XFILLER_46_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16923_ _14541_ VGND VGND VPWR VPWR _15413_ sky130_fd_sc_hd__buf_8
XFILLER_238_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29889_ registers\[18\]\[47\] _13033_ _13397_ VGND VGND VPWR VPWR _13405_ sky130_fd_sc_hd__mux2_1
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31920_ _14473_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19642_ _05095_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__clkbuf_8
XFILLER_238_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16854_ _15340_ _15345_ _15269_ VGND VGND VPWR VPWR _15346_ sky130_fd_sc_hd__o21ba_1
XFILLER_226_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19573_ registers\[56\]\[34\] registers\[57\]\[34\] registers\[58\]\[34\] registers\[59\]\[34\]
+ _06301_ _06091_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__mux4_1
XFILLER_18_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31851_ _14437_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16785_ _15273_ _15276_ _15277_ _15278_ VGND VGND VPWR VPWR _15279_ sky130_fd_sc_hd__o211a_1
XFILLER_19_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18524_ _05107_ _05281_ _05282_ _05117_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__a22o_1
X_30802_ _09756_ registers\[11\]\[31\] _13884_ VGND VGND VPWR VPWR _13886_ sky130_fd_sc_hd__mux2_1
XFILLER_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34570_ clknet_leaf_165_CLK _02684_ VGND VGND VPWR VPWR registers\[28\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31782_ registers\[59\]\[48\] net43 _14392_ VGND VGND VPWR VPWR _14401_ sky130_fd_sc_hd__mux2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33521_ clknet_leaf_361_CLK _01635_ VGND VGND VPWR VPWR registers\[44\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_30733_ registers\[12\]\[63\] _13066_ _13779_ VGND VGND VPWR VPWR _13849_ sky130_fd_sc_hd__mux2_1
XFILLER_179_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18455_ _05212_ _05215_ _05103_ _05105_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__o211a_1
XANTENNA_170 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17406_ _15684_ _15880_ _15881_ _15687_ VGND VGND VPWR VPWR _15882_ sky130_fd_sc_hd__a22o_1
XFILLER_159_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33452_ clknet_leaf_345_CLK _01566_ VGND VGND VPWR VPWR registers\[45\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18386_ _05058_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__buf_12
X_30664_ _13779_ VGND VGND VPWR VPWR _13813_ sky130_fd_sc_hd__buf_6
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32403_ clknet_leaf_104_CLK _00517_ VGND VGND VPWR VPWR registers\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36171_ clknet_leaf_164_CLK _04285_ VGND VGND VPWR VPWR registers\[49\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17337_ _15811_ _15814_ _15612_ VGND VGND VPWR VPWR _15815_ sky130_fd_sc_hd__o21ba_1
X_30595_ _13776_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33383_ clknet_leaf_59_CLK _01497_ VGND VGND VPWR VPWR registers\[46\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35122_ clknet_leaf_382_CLK _03236_ VGND VGND VPWR VPWR registers\[1\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_32334_ clknet_leaf_180_CLK _00448_ VGND VGND VPWR VPWR registers\[61\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17268_ registers\[44\]\[34\] registers\[45\]\[34\] registers\[46\]\[34\] registers\[47\]\[34\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15748_ sky130_fd_sc_hd__mux4_1
XFILLER_70_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19007_ registers\[48\]\[18\] registers\[49\]\[18\] registers\[50\]\[18\] registers\[51\]\[18\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__mux4_1
X_16219_ registers\[52\]\[4\] registers\[53\]\[4\] registers\[54\]\[4\] registers\[55\]\[4\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14729_ sky130_fd_sc_hd__mux4_1
X_35053_ clknet_leaf_395_CLK _03167_ VGND VGND VPWR VPWR registers\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_32265_ clknet_leaf_236_CLK _00379_ VGND VGND VPWR VPWR registers\[39\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17199_ registers\[32\]\[32\] registers\[33\]\[32\] registers\[34\]\[32\] registers\[35\]\[32\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15681_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_61_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_61_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34004_ clknet_leaf_119_CLK _02118_ VGND VGND VPWR VPWR registers\[36\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31216_ _14103_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32196_ clknet_leaf_399_CLK _00310_ VGND VGND VPWR VPWR registers\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31147_ _14067_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19909_ registers\[24\]\[43\] registers\[25\]\[43\] registers\[26\]\[43\] registers\[27\]\[43\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__mux4_1
Xclkbuf_6_29__f_CLK clknet_5_14_0_CLK VGND VGND VPWR VPWR clknet_6_29__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31078_ registers\[0\]\[34\] _13006_ _14026_ VGND VGND VPWR VPWR _14031_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35955_ clknet_leaf_380_CLK _04069_ VGND VGND VPWR VPWR registers\[6\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30029_ _13478_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__clkbuf_1
X_34906_ clknet_leaf_0_CLK _03020_ VGND VGND VPWR VPWR registers\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_22920_ net5 VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__buf_6
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35886_ clknet_leaf_391_CLK _04000_ VGND VGND VPWR VPWR registers\[7\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22851_ _09483_ _09486_ _07309_ VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__o21ba_1
X_34837_ clknet_leaf_96_CLK _02951_ VGND VGND VPWR VPWR registers\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21802_ _07324_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__clkbuf_4
X_25570_ _11011_ VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__buf_4
X_22782_ _09417_ _09420_ _07398_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__o21ba_1
X_34768_ clknet_leaf_111_CLK _02882_ VGND VGND VPWR VPWR registers\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24521_ _09590_ registers\[56\]\[36\] _10473_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__mux2_1
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21733_ registers\[60\]\[30\] registers\[61\]\[30\] registers\[62\]\[30\] registers\[63\]\[30\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__mux4_1
X_33719_ clknet_leaf_341_CLK _01833_ VGND VGND VPWR VPWR registers\[41\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34699_ clknet_leaf_149_CLK _02813_ VGND VGND VPWR VPWR registers\[26\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27240_ _11979_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24452_ _09521_ registers\[56\]\[3\] _10440_ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__mux2_1
X_21664_ _07328_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__buf_6
XFILLER_162_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23403_ registers\[39\]\[54\] _09806_ _09851_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27171_ _11943_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_990 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20615_ _07277_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__buf_12
X_24383_ registers\[57\]\[44\] _10397_ _10389_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__mux2_1
X_21595_ registers\[8\]\[26\] registers\[9\]\[26\] registers\[10\]\[26\] registers\[11\]\[26\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__mux4_1
XFILLER_197_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26122_ _10842_ registers\[45\]\[53\] _11356_ VGND VGND VPWR VPWR _11360_ sky130_fd_sc_hd__mux2_1
X_23334_ registers\[9\]\[59\] _09817_ _09798_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__mux2_1
X_20546_ registers\[32\]\[63\] registers\[33\]\[63\] registers\[34\]\[63\] registers\[35\]\[63\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__mux4_1
XFILLER_138_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26053_ _10772_ registers\[45\]\[20\] _11323_ VGND VGND VPWR VPWR _11324_ sky130_fd_sc_hd__mux2_1
XFILLER_192_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23265_ registers\[9\]\[38\] _09771_ _09754_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__mux2_1
XFILLER_106_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20477_ registers\[16\]\[60\] registers\[17\]\[60\] registers\[18\]\[60\] registers\[19\]\[60\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__mux4_1
XFILLER_119_994 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_52_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25004_ net45 VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__buf_4
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22216_ _08848_ _08855_ _08864_ _08871_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__or4_4
XFILLER_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23196_ _09728_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29812_ registers\[18\]\[10\] _12955_ _13364_ VGND VGND VPWR VPWR _13365_ sky130_fd_sc_hd__mux2_1
XANTENNA_1508 _07395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22147_ _08804_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_2
XTAP_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1519 _08841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29743_ _13328_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__clkbuf_1
X_26955_ _11819_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__clkbuf_1
X_22078_ registers\[44\]\[40\] registers\[45\]\[40\] registers\[46\]\[40\] registers\[47\]\[40\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__mux4_1
XTAP_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21029_ _07648_ _07716_ _07717_ _07652_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__a22o_1
X_25906_ _11246_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29674_ registers\[1\]\[9\] _12953_ _13282_ VGND VGND VPWR VPWR _13292_ sky130_fd_sc_hd__mux2_1
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26886_ _11771_ registers\[3\]\[20\] _11772_ VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__mux2_1
XFILLER_87_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28625_ _11845_ registers\[27\]\[55\] _12703_ VGND VGND VPWR VPWR _12709_ sky130_fd_sc_hd__mux2_1
X_25837_ _10827_ registers\[47\]\[46\] _11203_ VGND VGND VPWR VPWR _11210_ sky130_fd_sc_hd__mux2_1
XFILLER_207_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28556_ _11776_ registers\[27\]\[22\] _12670_ VGND VGND VPWR VPWR _12673_ sky130_fd_sc_hd__mux2_1
X_16570_ _14541_ VGND VGND VPWR VPWR _15070_ sky130_fd_sc_hd__clkbuf_8
X_25768_ _10758_ registers\[47\]\[13\] _11170_ VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__mux2_1
XFILLER_28_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27507_ _11809_ registers\[35\]\[38\] _12111_ VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__mux2_1
X_24719_ _10512_ _10585_ VGND VGND VPWR VPWR _10586_ sky130_fd_sc_hd__nand2_8
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28487_ _12636_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__clkbuf_1
X_25699_ _11136_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18240_ registers\[20\]\[62\] registers\[21\]\[62\] registers\[22\]\[62\] registers\[23\]\[62\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__mux4_1
XFILLER_163_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27438_ _11740_ registers\[35\]\[5\] _12078_ VGND VGND VPWR VPWR _12084_ sky130_fd_sc_hd__mux2_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18171_ _14491_ _04936_ _04937_ _14501_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__a22o_1
XFILLER_129_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27369_ _12047_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29108_ registers\[23\]\[18\] _12972_ _12956_ VGND VGND VPWR VPWR _12973_ sky130_fd_sc_hd__mux2_1
X_17122_ _15334_ _15604_ _15605_ _15339_ VGND VGND VPWR VPWR _15606_ sky130_fd_sc_hd__a22o_1
XFILLER_129_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30380_ _09730_ registers\[14\]\[23\] _13660_ VGND VGND VPWR VPWR _13664_ sky130_fd_sc_hd__mux2_1
XFILLER_128_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17053_ _15341_ _15537_ _15538_ _15344_ VGND VGND VPWR VPWR _15539_ sky130_fd_sc_hd__a22o_1
X_29039_ _12926_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_43_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_43_CLK sky130_fd_sc_hd__clkbuf_16
X_16004_ _14492_ VGND VGND VPWR VPWR _14518_ sky130_fd_sc_hd__buf_12
XFILLER_87_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32050_ clknet_leaf_380_CLK _00228_ VGND VGND VPWR VPWR registers\[62\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31001_ registers\[10\]\[62\] _13064_ _13921_ VGND VGND VPWR VPWR _13990_ sky130_fd_sc_hd__mux2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17955_ _04481_ _04727_ _04728_ _04484_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__a22o_1
XFILLER_140_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16906_ registers\[28\]\[23\] registers\[29\]\[23\] registers\[30\]\[23\] registers\[31\]\[23\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15397_ sky130_fd_sc_hd__mux4_1
X_35740_ clknet_leaf_478_CLK _03854_ VGND VGND VPWR VPWR registers\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32952_ clknet_leaf_331_CLK _01066_ VGND VGND VPWR VPWR registers\[53\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17886_ registers\[0\]\[51\] registers\[1\]\[51\] registers\[2\]\[51\] registers\[3\]\[51\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__mux4_1
X_19625_ registers\[28\]\[35\] registers\[29\]\[35\] registers\[30\]\[35\] registers\[31\]\[35\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__mux4_1
XFILLER_93_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31903_ _09778_ registers\[49\]\[41\] _14463_ VGND VGND VPWR VPWR _14465_ sky130_fd_sc_hd__mux2_1
X_35671_ clknet_leaf_85_CLK _03785_ VGND VGND VPWR VPWR registers\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_16837_ registers\[20\]\[21\] registers\[21\]\[21\] registers\[22\]\[21\] registers\[23\]\[21\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15330_ sky130_fd_sc_hd__mux4_1
X_32883_ clknet_leaf_355_CLK _00997_ VGND VGND VPWR VPWR registers\[54\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34622_ clknet_leaf_179_CLK _02736_ VGND VGND VPWR VPWR registers\[27\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31834_ _14428_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__clkbuf_1
X_19556_ registers\[24\]\[33\] registers\[25\]\[33\] registers\[26\]\[33\] registers\[27\]\[33\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__mux4_1
Xclkbuf_5_22_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_22_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16768_ registers\[32\]\[20\] registers\[33\]\[20\] registers\[34\]\[20\] registers\[35\]\[20\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15262_ sky130_fd_sc_hd__mux4_1
XFILLER_185_1250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18507_ registers\[32\]\[4\] registers\[33\]\[4\] registers\[34\]\[4\] registers\[35\]\[4\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__mux4_1
XFILLER_206_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34553_ clknet_leaf_185_CLK _02667_ VGND VGND VPWR VPWR registers\[28\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31765_ _14347_ VGND VGND VPWR VPWR _14392_ sky130_fd_sc_hd__buf_4
X_19487_ registers\[16\]\[31\] registers\[17\]\[31\] registers\[18\]\[31\] registers\[19\]\[31\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__mux4_1
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16699_ registers\[36\]\[18\] registers\[37\]\[18\] registers\[38\]\[18\] registers\[39\]\[18\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15195_ sky130_fd_sc_hd__mux4_1
X_33504_ clknet_leaf_34_CLK _01618_ VGND VGND VPWR VPWR registers\[44\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_30716_ _13840_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__clkbuf_1
X_18438_ _05045_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__buf_6
XFILLER_142_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34484_ clknet_leaf_414_CLK _02598_ VGND VGND VPWR VPWR registers\[2\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31696_ registers\[59\]\[7\] net62 _14348_ VGND VGND VPWR VPWR _14356_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36223_ clknet_leaf_117_CLK _00107_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dfxtp_1
X_33435_ clknet_leaf_31_CLK _01549_ VGND VGND VPWR VPWR registers\[45\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18369_ _05119_ _05124_ _05129_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__a22o_1
X_30647_ _13804_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__clkbuf_1
X_20400_ _06919_ _07103_ _07104_ _06922_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__a22o_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36154_ clknet_leaf_281_CLK _04268_ VGND VGND VPWR VPWR registers\[49\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_33366_ clknet_leaf_122_CLK _01480_ VGND VGND VPWR VPWR registers\[46\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21380_ registers\[60\]\[20\] registers\[61\]\[20\] registers\[62\]\[20\] registers\[63\]\[20\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__mux4_1
X_30578_ _09804_ registers\[13\]\[53\] _13764_ VGND VGND VPWR VPWR _13768_ sky130_fd_sc_hd__mux2_1
XFILLER_120_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35105_ clknet_leaf_488_CLK _03219_ VGND VGND VPWR VPWR registers\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_20331_ _06873_ _07037_ _07038_ _06878_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__a22o_1
XFILLER_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32317_ clknet_leaf_191_CLK _00431_ VGND VGND VPWR VPWR registers\[19\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36085_ clknet_leaf_351_CLK _04199_ VGND VGND VPWR VPWR registers\[59\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_33297_ clknet_leaf_129_CLK _01411_ VGND VGND VPWR VPWR registers\[47\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_34_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_34_CLK sky130_fd_sc_hd__clkbuf_16
X_23050_ net51 VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35036_ clknet_leaf_491_CLK _03150_ VGND VGND VPWR VPWR registers\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_20262_ registers\[24\]\[53\] registers\[25\]\[53\] registers\[26\]\[53\] registers\[27\]\[53\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__mux4_1
XFILLER_227_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32248_ clknet_leaf_337_CLK _00362_ VGND VGND VPWR VPWR registers\[39\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22001_ registers\[40\]\[38\] registers\[41\]\[38\] registers\[42\]\[38\] registers\[43\]\[38\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__mux4_1
XTAP_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20193_ registers\[16\]\[51\] registers\[17\]\[51\] registers\[18\]\[51\] registers\[19\]\[51\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__mux4_1
XFILLER_66_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32179_ clknet_leaf_15_CLK _00293_ VGND VGND VPWR VPWR registers\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23952_ _09628_ registers\[60\]\[54\] _10144_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__mux2_1
XFILLER_130_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26740_ registers\[40\]\[25\] _10357_ _11680_ VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__mux2_1
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35938_ clknet_leaf_469_CLK _04052_ VGND VGND VPWR VPWR registers\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22903_ _09530_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26671_ _10850_ registers\[41\]\[57\] _11641_ VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__mux2_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35869_ clknet_leaf_476_CLK _03983_ VGND VGND VPWR VPWR registers\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_23883_ _09559_ registers\[60\]\[21\] _10111_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__mux2_1
XFILLER_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_906 _09676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28410_ _11765_ registers\[28\]\[17\] _12588_ VGND VGND VPWR VPWR _12596_ sky130_fd_sc_hd__mux2_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1088 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22834_ _07296_ _09469_ _09470_ _07302_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__a22o_1
X_25622_ registers\[48\]\[9\] _10323_ _11086_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__mux2_1
X_29390_ _09662_ registers\[21\]\[2\] _13140_ VGND VGND VPWR VPWR _13143_ sky130_fd_sc_hd__mux2_1
XANTENNA_917 _09758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_928 _09869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_939 _10288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28341_ _12559_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__clkbuf_1
X_25553_ _11058_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__clkbuf_1
X_22765_ registers\[60\]\[60\] registers\[61\]\[60\] registers\[62\]\[60\] registers\[63\]\[60\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__mux4_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24504_ _09573_ registers\[56\]\[28\] _10462_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21716_ _08080_ _08384_ _08385_ _08085_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__a22o_1
X_28272_ _12523_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25484_ registers\[4\]\[9\] _10323_ _11012_ VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22696_ registers\[32\]\[58\] registers\[33\]\[58\] registers\[34\]\[58\] registers\[35\]\[58\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__mux4_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24435_ registers\[57\]\[61\] _10432_ net283 VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__mux2_1
XFILLER_169_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27223_ _11795_ registers\[37\]\[31\] _11969_ VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__mux2_1
X_21647_ _08318_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27154_ _11861_ registers\[38\]\[63\] _11864_ VGND VGND VPWR VPWR _11934_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24366_ net33 VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__buf_4
XANTENNA_70 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21578_ registers\[40\]\[26\] registers\[41\]\[26\] registers\[42\]\[26\] registers\[43\]\[26\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__mux4_1
XANTENNA_81 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26105_ _10825_ registers\[45\]\[45\] _11345_ VGND VGND VPWR VPWR _11351_ sky130_fd_sc_hd__mux2_1
X_23317_ registers\[9\]\[54\] _09806_ _09798_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__mux2_1
XANTENNA_92 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20529_ registers\[8\]\[62\] registers\[9\]\[62\] registers\[10\]\[62\] registers\[11\]\[62\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__mux4_1
XFILLER_153_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27085_ _11864_ VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__buf_4
XFILLER_153_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24297_ _10339_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_25_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_25_CLK sky130_fd_sc_hd__clkbuf_16
X_26036_ _10756_ registers\[45\]\[12\] _11312_ VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__mux2_1
X_23248_ registers\[9\]\[33\] _09760_ _09754_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23179_ _09719_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
XTAP_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1305 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1316 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1327 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1338 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27987_ _12373_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1349 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _04481_ _04518_ _04519_ _04484_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__a22o_1
X_29726_ _13319_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26938_ _11807_ registers\[3\]\[37\] _11793_ VGND VGND VPWR VPWR _11808_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_12__f_CLK clknet_5_6_0_CLK VGND VGND VPWR VPWR clknet_6_12__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29657_ _13283_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__clkbuf_1
X_17671_ registers\[12\]\[45\] registers\[13\]\[45\] registers\[14\]\[45\] registers\[15\]\[45\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__mux4_1
XFILLER_101_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26869_ net7 VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__buf_4
X_19410_ _06140_ _06143_ _05837_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__o21ba_1
XFILLER_1_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28608_ _11828_ registers\[27\]\[47\] _12692_ VGND VGND VPWR VPWR _12700_ sky130_fd_sc_hd__mux2_1
X_16622_ _15117_ _15120_ _14959_ VGND VGND VPWR VPWR _15121_ sky130_fd_sc_hd__o21ba_1
XFILLER_235_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_235_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29588_ registers\[20\]\[32\] _13002_ _13244_ VGND VGND VPWR VPWR _13247_ sky130_fd_sc_hd__mux2_1
XFILLER_28_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _05839_ _06075_ _06076_ _05842_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a22o_1
X_16553_ registers\[28\]\[13\] registers\[29\]\[13\] registers\[30\]\[13\] registers\[31\]\[13\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15054_ sky130_fd_sc_hd__mux4_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28539_ _11759_ registers\[27\]\[14\] _12659_ VGND VGND VPWR VPWR _12664_ sky130_fd_sc_hd__mux2_1
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31550_ _14279_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19272_ registers\[28\]\[25\] registers\[29\]\[25\] registers\[30\]\[25\] registers\[31\]\[25\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16484_ registers\[20\]\[11\] registers\[21\]\[11\] registers\[22\]\[11\] registers\[23\]\[11\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _14987_ sky130_fd_sc_hd__mux4_1
X_18223_ registers\[48\]\[62\] registers\[49\]\[62\] registers\[50\]\[62\] registers\[51\]\[62\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__mux4_1
X_30501_ _13727_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31481_ _09760_ registers\[6\]\[33\] _14239_ VGND VGND VPWR VPWR _14243_ sky130_fd_sc_hd__mux2_1
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33220_ clknet_leaf_231_CLK _01334_ VGND VGND VPWR VPWR registers\[4\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18154_ _04921_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_2
XFILLER_175_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30432_ _09793_ registers\[14\]\[48\] _13682_ VGND VGND VPWR VPWR _13691_ sky130_fd_sc_hd__mux2_1
XFILLER_129_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17105_ registers\[0\]\[29\] registers\[1\]\[29\] registers\[2\]\[29\] registers\[3\]\[29\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15590_ sky130_fd_sc_hd__mux4_1
X_33151_ clknet_leaf_268_CLK _01265_ VGND VGND VPWR VPWR registers\[50\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18085_ _04851_ _04854_ _04630_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__o21ba_1
X_30363_ _09689_ registers\[14\]\[15\] _13649_ VGND VGND VPWR VPWR _13655_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_16_CLK sky130_fd_sc_hd__clkbuf_16
X_32102_ clknet_leaf_483_CLK _00016_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dfxtp_1
X_17036_ registers\[4\]\[27\] registers\[5\]\[27\] registers\[6\]\[27\] registers\[7\]\[27\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15523_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30294_ registers\[15\]\[47\] _13033_ _13610_ VGND VGND VPWR VPWR _13618_ sky130_fd_sc_hd__mux2_1
X_33082_ clknet_leaf_281_CLK _01196_ VGND VGND VPWR VPWR registers\[51\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_32033_ clknet_leaf_444_CLK _00211_ VGND VGND VPWR VPWR registers\[62\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ registers\[16\]\[17\] registers\[17\]\[17\] registers\[18\]\[17\] registers\[19\]\[17\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__mux4_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17938_ _04712_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_2
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33984_ clknet_leaf_260_CLK _02098_ VGND VGND VPWR VPWR registers\[37\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35723_ clknet_leaf_151_CLK _03837_ VGND VGND VPWR VPWR registers\[10\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32935_ clknet_leaf_437_CLK _01049_ VGND VGND VPWR VPWR registers\[53\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17869_ _04612_ _04621_ _04631_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__or4_4
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19608_ _06090_ _06334_ _06335_ _06096_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__a22o_1
X_35654_ clknet_leaf_215_CLK _03768_ VGND VGND VPWR VPWR registers\[11\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20880_ registers\[48\]\[6\] registers\[49\]\[6\] registers\[50\]\[6\] registers\[51\]\[6\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__mux4_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32866_ clknet_leaf_444_CLK _00980_ VGND VGND VPWR VPWR registers\[54\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34605_ clknet_leaf_403_CLK _02719_ VGND VGND VPWR VPWR registers\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31817_ _09648_ registers\[49\]\[0\] _14419_ VGND VGND VPWR VPWR _14420_ sky130_fd_sc_hd__mux2_1
X_19539_ _06265_ _06268_ _06161_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35585_ clknet_leaf_236_CLK _03699_ VGND VGND VPWR VPWR registers\[12\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32797_ clknet_leaf_55_CLK _00911_ VGND VGND VPWR VPWR registers\[55\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_22550_ registers\[52\]\[53\] registers\[53\]\[53\] registers\[54\]\[53\] registers\[55\]\[53\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__mux4_1
X_34536_ clknet_leaf_453_CLK _02650_ VGND VGND VPWR VPWR registers\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31748_ _14383_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21501_ _07929_ _08175_ _08176_ _07932_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__a22o_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22481_ registers\[60\]\[51\] registers\[61\]\[51\] registers\[62\]\[51\] registers\[63\]\[51\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__mux4_1
X_34467_ clknet_leaf_471_CLK _02581_ VGND VGND VPWR VPWR registers\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31679_ _14346_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24220_ _09624_ registers\[58\]\[52\] _10288_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__mux2_1
X_36206_ clknet_leaf_100_CLK _00089_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dfxtp_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33418_ clknet_leaf_163_CLK _01532_ VGND VGND VPWR VPWR registers\[46\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_21432_ _08106_ _08109_ _08073_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__o21ba_1
XFILLER_124_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34398_ clknet_leaf_492_CLK _02512_ VGND VGND VPWR VPWR registers\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24151_ _10254_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__clkbuf_1
X_36137_ clknet_leaf_424_CLK _04251_ VGND VGND VPWR VPWR registers\[49\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_33349_ clknet_leaf_256_CLK _01463_ VGND VGND VPWR VPWR registers\[47\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_21363_ _07737_ _08041_ _08042_ _07742_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__a22o_1
XFILLER_175_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23102_ net56 VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__buf_4
X_20314_ _06776_ _07020_ _07021_ _06782_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__a22o_1
X_24082_ _09622_ registers\[5\]\[51\] _10216_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__mux2_1
XFILLER_163_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36068_ clknet_leaf_441_CLK _04182_ VGND VGND VPWR VPWR registers\[59\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_21294_ _07975_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35019_ clknet_leaf_143_CLK _03133_ VGND VGND VPWR VPWR registers\[21\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_23033_ _09618_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
X_27910_ registers\[32\]\[36\] _10380_ _12326_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__mux2_1
XFILLER_239_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20245_ _06951_ _06954_ _06847_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__o21ba_1
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28890_ _12848_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27841_ registers\[32\]\[3\] _10311_ _12293_ VGND VGND VPWR VPWR _12297_ sky130_fd_sc_hd__mux2_1
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20176_ _06576_ _06886_ _06887_ _06579_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__a22o_1
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27772_ _12260_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__clkbuf_1
X_24984_ _10725_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__clkbuf_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29511_ _09819_ registers\[21\]\[60\] _13139_ VGND VGND VPWR VPWR _13206_ sky130_fd_sc_hd__mux2_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26723_ registers\[40\]\[17\] _10340_ _11669_ VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__mux2_1
XFILLER_217_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _09611_ registers\[60\]\[46\] _10133_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__mux2_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29442_ _09747_ registers\[21\]\[27\] _13162_ VGND VGND VPWR VPWR _13170_ sky130_fd_sc_hd__mux2_1
X_26654_ _10833_ registers\[41\]\[49\] _11630_ VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__mux2_1
XFILLER_131_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23866_ _09542_ registers\[60\]\[13\] _10100_ VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__mux2_1
XANTENNA_703 _07281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_714 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_725 _07349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_736 _07356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22817_ _07313_ _09452_ _09453_ _07322_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__a22o_1
X_25605_ _11087_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_747 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29373_ _13133_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23797_ _09609_ registers\[29\]\[45\] _10061_ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__mux2_1
XANTENNA_758 _07392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26585_ _10764_ registers\[41\]\[16\] _11597_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_769 _07802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28324_ registers\[2\]\[40\] _10388_ _12550_ VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__mux2_1
X_22748_ _09104_ _09386_ _09387_ _09107_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__a22o_1
X_25536_ _11049_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25467_ _11013_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_1
X_28255_ _12514_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__clkbuf_1
X_22679_ registers\[8\]\[57\] registers\[9\]\[57\] registers\[10\]\[57\] registers\[11\]\[57\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__mux4_1
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24418_ _10421_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27206_ _11778_ registers\[37\]\[23\] _11958_ VGND VGND VPWR VPWR _11962_ sky130_fd_sc_hd__mux2_1
XFILLER_173_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25398_ _10802_ registers\[50\]\[34\] _10970_ VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__mux2_1
X_28186_ _11811_ registers\[30\]\[39\] _12468_ VGND VGND VPWR VPWR _12478_ sky130_fd_sc_hd__mux2_1
XFILLER_126_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27137_ _11925_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_1
X_24349_ registers\[57\]\[33\] _10374_ _10368_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__mux2_1
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27068_ _11889_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26019_ _10739_ registers\[45\]\[4\] _11301_ VGND VGND VPWR VPWR _11306_ sky130_fd_sc_hd__mux2_1
XFILLER_180_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18910_ registers\[0\]\[15\] registers\[1\]\[15\] registers\[2\]\[15\] registers\[3\]\[15\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__mux4_1
XTAP_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19890_ registers\[36\]\[43\] registers\[37\]\[43\] registers\[38\]\[43\] registers\[39\]\[43\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__mux4_1
XFILLER_10_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1102 _14539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1113 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18841_ registers\[8\]\[13\] registers\[9\]\[13\] registers\[10\]\[13\] registers\[11\]\[13\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__mux4_1
XTAP_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1124 _14584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1135 _14613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1146 _15547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1157 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18772_ _05520_ _05523_ _05483_ _05484_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o211a_2
XFILLER_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1168 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15984_ registers\[40\]\[0\] registers\[41\]\[0\] registers\[42\]\[0\] registers\[43\]\[0\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _14498_ sky130_fd_sc_hd__mux4_1
XTAP_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1179 _15777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17723_ registers\[32\]\[47\] registers\[33\]\[47\] registers\[34\]\[47\] registers\[35\]\[47\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__mux4_1
X_29709_ _13310_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__clkbuf_1
XTAP_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30981_ registers\[10\]\[52\] _13044_ _13977_ VGND VGND VPWR VPWR _13980_ sky130_fd_sc_hd__mux2_1
XTAP_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32720_ clknet_leaf_173_CLK _00834_ VGND VGND VPWR VPWR registers\[56\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17654_ _04333_ _04434_ _04435_ _04338_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__a22o_1
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_5_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16605_ _14863_ _15102_ _15103_ _14867_ VGND VGND VPWR VPWR _15104_ sky130_fd_sc_hd__a22o_1
X_32651_ clknet_leaf_164_CLK _00765_ VGND VGND VPWR VPWR registers\[58\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_17585_ _04369_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31602_ _14306_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__clkbuf_1
X_19324_ _06054_ _06059_ _05818_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__o21ba_1
X_16536_ _14855_ _15035_ _15036_ _14861_ VGND VGND VPWR VPWR _15037_ sky130_fd_sc_hd__a22o_1
X_35370_ clknet_leaf_398_CLK _03484_ VGND VGND VPWR VPWR registers\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_32582_ clknet_leaf_210_CLK _00696_ VGND VGND VPWR VPWR registers\[5\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34321_ clknet_leaf_101_CLK _02435_ VGND VGND VPWR VPWR registers\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31533_ _09815_ registers\[6\]\[58\] _14261_ VGND VGND VPWR VPWR _14270_ sky130_fd_sc_hd__mux2_1
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19255_ _05747_ _05991_ _05992_ _05753_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__a22o_1
XFILLER_177_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16467_ registers\[48\]\[11\] registers\[49\]\[11\] registers\[50\]\[11\] registers\[51\]\[11\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _14970_ sky130_fd_sc_hd__mux4_1
XFILLER_176_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18206_ registers\[24\]\[61\] registers\[25\]\[61\] registers\[26\]\[61\] registers\[27\]\[61\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__mux4_1
X_34252_ clknet_leaf_168_CLK _02366_ VGND VGND VPWR VPWR registers\[33\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_31464_ _09742_ registers\[6\]\[25\] _14228_ VGND VGND VPWR VPWR _14234_ sky130_fd_sc_hd__mux2_1
X_19186_ _05922_ _05925_ _05818_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__o21ba_1
X_16398_ registers\[8\]\[9\] registers\[9\]\[9\] registers\[10\]\[9\] registers\[11\]\[9\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14903_ sky130_fd_sc_hd__mux4_1
XFILLER_30_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33203_ clknet_leaf_380_CLK _01317_ VGND VGND VPWR VPWR registers\[4\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_18137_ _14600_ _04903_ _04904_ _14610_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__a22o_1
XFILLER_145_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30415_ _13637_ VGND VGND VPWR VPWR _13682_ sky130_fd_sc_hd__buf_4
X_34183_ clknet_leaf_244_CLK _02297_ VGND VGND VPWR VPWR registers\[34\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_31395_ _14197_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33134_ clknet_leaf_372_CLK _01248_ VGND VGND VPWR VPWR registers\[50\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_18068_ registers\[44\]\[57\] registers\[45\]\[57\] registers\[46\]\[57\] registers\[47\]\[57\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__mux4_1
X_30346_ _09672_ registers\[14\]\[7\] _13638_ VGND VGND VPWR VPWR _13646_ sky130_fd_sc_hd__mux2_1
XFILLER_144_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17019_ registers\[44\]\[27\] registers\[45\]\[27\] registers\[46\]\[27\] registers\[47\]\[27\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15506_ sky130_fd_sc_hd__mux4_1
XFILLER_154_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33065_ clknet_leaf_435_CLK _01179_ VGND VGND VPWR VPWR registers\[51\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30277_ registers\[15\]\[39\] _13016_ _13599_ VGND VGND VPWR VPWR _13609_ sky130_fd_sc_hd__mux2_1
X_32016_ clknet_leaf_175_CLK _00194_ VGND VGND VPWR VPWR registers\[62\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_20030_ _06740_ _06745_ _06504_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__o21ba_1
XFILLER_67_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1680 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1691 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21981_ registers\[60\]\[37\] registers\[61\]\[37\] registers\[62\]\[37\] registers\[63\]\[37\]
+ _08541_ _08335_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__mux4_1
X_33967_ clknet_leaf_356_CLK _02081_ VGND VGND VPWR VPWR registers\[37\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23720_ _10026_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20932_ _07620_ _07623_ _07370_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__o21ba_1
X_32918_ clknet_leaf_62_CLK _01032_ VGND VGND VPWR VPWR registers\[53\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35706_ clknet_leaf_302_CLK _03820_ VGND VGND VPWR VPWR registers\[10\]\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33898_ clknet_leaf_427_CLK _02012_ VGND VGND VPWR VPWR registers\[38\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23651_ registers\[61\]\[41\] _09778_ _09987_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__mux2_1
X_32849_ clknet_leaf_173_CLK _00963_ VGND VGND VPWR VPWR registers\[54\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_20863_ registers\[24\]\[5\] registers\[25\]\[5\] registers\[26\]\[5\] registers\[27\]\[5\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__mux4_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35637_ clknet_leaf_324_CLK _03751_ VGND VGND VPWR VPWR registers\[11\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22602_ _09243_ _09246_ _09116_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__o21ba_1
XFILLER_228_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26370_ _11490_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23582_ _09952_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
X_35568_ clknet_leaf_375_CLK _03682_ VGND VGND VPWR VPWR registers\[12\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_20794_ registers\[4\]\[3\] registers\[5\]\[3\] registers\[6\]\[3\] registers\[7\]\[3\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__mux4_1
XFILLER_74_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25321_ _10933_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__clkbuf_1
X_22533_ registers\[28\]\[52\] registers\[29\]\[52\] registers\[30\]\[52\] registers\[31\]\[52\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__mux4_1
X_34519_ clknet_leaf_98_CLK _02633_ VGND VGND VPWR VPWR registers\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_35499_ clknet_leaf_397_CLK _03613_ VGND VGND VPWR VPWR registers\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28040_ _12401_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__clkbuf_1
X_25252_ _10897_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_1
X_22464_ registers\[20\]\[50\] registers\[21\]\[50\] registers\[22\]\[50\] registers\[23\]\[50\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__mux4_1
XFILLER_183_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24203_ _09607_ registers\[58\]\[44\] _10277_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__mux2_1
X_21415_ registers\[44\]\[21\] registers\[45\]\[21\] registers\[46\]\[21\] registers\[47\]\[21\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__mux4_1
X_25183_ net59 VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__buf_2
X_22395_ _07287_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__clkbuf_8
XFILLER_202_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24134_ _09538_ registers\[58\]\[11\] _10244_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__mux2_1
XFILLER_108_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21346_ _07983_ _08024_ _08025_ _07989_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__a22o_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29991_ registers\[17\]\[31\] _13000_ _13457_ VGND VGND VPWR VPWR _13459_ sky130_fd_sc_hd__mux2_1
XFILLER_190_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24065_ _09605_ registers\[5\]\[43\] _10205_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__mux2_1
X_28942_ registers\[24\]\[13\] _10332_ _12872_ VGND VGND VPWR VPWR _12876_ sky130_fd_sc_hd__mux2_1
XFILLER_235_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21277_ _07648_ _07957_ _07958_ _07652_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__a22o_1
XFILLER_172_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23016_ net39 VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20228_ registers\[24\]\[52\] registers\[25\]\[52\] registers\[26\]\[52\] registers\[27\]\[52\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__mux4_1
XFILLER_235_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28873_ _12839_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27824_ _12287_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__clkbuf_1
X_20159_ _06868_ _06869_ _06870_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__a22o_1
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27755_ _12251_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__clkbuf_1
X_24967_ _09626_ registers\[53\]\[53\] _10713_ VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__mux2_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26706_ registers\[40\]\[9\] _10323_ _11658_ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__mux2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23918_ _09594_ registers\[60\]\[38\] _10122_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__mux2_1
X_27686_ registers\[34\]\[58\] _10426_ _12206_ VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__mux2_1
XFILLER_206_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_500 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24898_ _09556_ registers\[53\]\[20\] _10680_ VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__mux2_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_511 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29425_ _09697_ registers\[21\]\[19\] _13151_ VGND VGND VPWR VPWR _13161_ sky130_fd_sc_hd__mux2_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_522 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_533 _00176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26637_ _11631_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__clkbuf_1
X_23849_ _09525_ registers\[60\]\[5\] _10089_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__mux2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_544 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_555 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_566 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_577 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29356_ _09797_ registers\[22\]\[50\] _13124_ VGND VGND VPWR VPWR _13125_ sky130_fd_sc_hd__mux2_1
X_17370_ registers\[32\]\[37\] registers\[33\]\[37\] registers\[34\]\[37\] registers\[35\]\[37\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15847_ sky130_fd_sc_hd__mux4_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26568_ _10747_ registers\[41\]\[8\] _11586_ VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__mux2_1
XANTENNA_588 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_599 _05088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16321_ _14528_ _14826_ _14827_ _14537_ VGND VGND VPWR VPWR _14828_ sky130_fd_sc_hd__a22o_1
X_28307_ registers\[2\]\[32\] _10372_ _12539_ VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__mux2_1
XFILLER_14_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25519_ _11040_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29287_ _13088_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__clkbuf_1
X_26499_ _11513_ VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__buf_4
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19040_ registers\[44\]\[19\] registers\[45\]\[19\] registers\[46\]\[19\] registers\[47\]\[19\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__mux4_1
X_28238_ _11008_ _12149_ VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__nor2_8
XFILLER_220_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16252_ _14540_ _14759_ _14760_ _14551_ VGND VGND VPWR VPWR _14761_ sky130_fd_sc_hd__a22o_1
XFILLER_103_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16183_ _14528_ _14692_ _14693_ _14537_ VGND VGND VPWR VPWR _14694_ sky130_fd_sc_hd__a22o_1
X_28169_ _12469_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__clkbuf_1
X_30200_ registers\[15\]\[2\] _12939_ _13566_ VGND VGND VPWR VPWR _13569_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput209 net209 VGND VGND VPWR VPWR D2[5] sky130_fd_sc_hd__buf_2
X_31180_ _14084_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19942_ _05113_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__buf_6
X_30131_ _13532_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30062_ _13496_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19873_ _06379_ _06592_ _06593_ _06382_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__a22o_1
XFILLER_218_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18824_ _05569_ _05574_ _05508_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__o21ba_1
XFILLER_96_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34870_ clknet_leaf_308_CLK _02984_ VGND VGND VPWR VPWR registers\[23\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33821_ clknet_leaf_478_CLK _01935_ VGND VGND VPWR VPWR registers\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _05162_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__buf_2
XFILLER_62_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17706_ registers\[12\]\[46\] registers\[13\]\[46\] registers\[14\]\[46\] registers\[15\]\[46\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__mux4_1
XFILLER_188_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33752_ clknet_leaf_86_CLK _01866_ VGND VGND VPWR VPWR registers\[40\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_18686_ _05197_ _05436_ _05439_ _05202_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__a22o_1
XFILLER_149_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30964_ registers\[10\]\[44\] _13027_ _13966_ VGND VGND VPWR VPWR _13971_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32703_ clknet_leaf_290_CLK _00817_ VGND VGND VPWR VPWR registers\[57\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17637_ registers\[12\]\[44\] registers\[13\]\[44\] registers\[14\]\[44\] registers\[15\]\[44\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__mux4_1
X_33683_ clknet_leaf_127_CLK _01797_ VGND VGND VPWR VPWR registers\[41\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30895_ registers\[10\]\[11\] _12958_ _13933_ VGND VGND VPWR VPWR _13935_ sky130_fd_sc_hd__mux2_1
X_35422_ clknet_leaf_483_CLK _03536_ VGND VGND VPWR VPWR registers\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_32634_ clknet_leaf_286_CLK _00748_ VGND VGND VPWR VPWR registers\[58\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_17568_ registers\[8\]\[42\] registers\[9\]\[42\] registers\[10\]\[42\] registers\[11\]\[42\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__mux4_1
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19307_ _05143_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__buf_4
XFILLER_56_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16519_ _14592_ VGND VGND VPWR VPWR _15021_ sky130_fd_sc_hd__buf_6
XFILLER_56_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35353_ clknet_leaf_13_CLK _03467_ VGND VGND VPWR VPWR registers\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_32565_ clknet_leaf_323_CLK _00679_ VGND VGND VPWR VPWR registers\[5\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_17499_ _15830_ _15971_ _15972_ _15833_ VGND VGND VPWR VPWR _15973_ sky130_fd_sc_hd__a22o_1
XFILLER_225_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34304_ clknet_leaf_258_CLK _02418_ VGND VGND VPWR VPWR registers\[32\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_31516_ _14205_ VGND VGND VPWR VPWR _14261_ sky130_fd_sc_hd__buf_4
XFILLER_177_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19238_ registers\[16\]\[24\] registers\[17\]\[24\] registers\[18\]\[24\] registers\[19\]\[24\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__mux4_1
X_35284_ clknet_leaf_93_CLK _03398_ VGND VGND VPWR VPWR registers\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32496_ clknet_leaf_368_CLK _00610_ VGND VGND VPWR VPWR registers\[60\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34235_ clknet_leaf_279_CLK _02349_ VGND VGND VPWR VPWR registers\[33\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31447_ _09693_ registers\[6\]\[17\] _14217_ VGND VGND VPWR VPWR _14225_ sky130_fd_sc_hd__mux2_1
X_19169_ registers\[24\]\[22\] registers\[25\]\[22\] registers\[26\]\[22\] registers\[27\]\[22\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__mux4_1
XFILLER_30_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21200_ registers\[56\]\[15\] registers\[57\]\[15\] registers\[58\]\[15\] registers\[59\]\[15\]
+ _07851_ _07641_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__mux4_1
X_22180_ registers\[28\]\[42\] registers\[29\]\[42\] registers\[30\]\[42\] registers\[31\]\[42\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34166_ clknet_leaf_342_CLK _02280_ VGND VGND VPWR VPWR registers\[34\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_31378_ _14188_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33117_ clknet_leaf_51_CLK _01231_ VGND VGND VPWR VPWR registers\[50\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_21131_ registers\[36\]\[13\] registers\[37\]\[13\] registers\[38\]\[13\] registers\[39\]\[13\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__mux4_1
X_30329_ _09651_ _09649_ _09650_ VGND VGND VPWR VPWR _13636_ sky130_fd_sc_hd__nor3b_4
XFILLER_160_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34097_ clknet_leaf_355_CLK _02211_ VGND VGND VPWR VPWR registers\[35\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33048_ clknet_leaf_52_CLK _01162_ VGND VGND VPWR VPWR registers\[51\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_21062_ registers\[44\]\[11\] registers\[45\]\[11\] registers\[46\]\[11\] registers\[47\]\[11\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__mux4_1
XFILLER_236_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20013_ _05081_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__buf_4
XFILLER_141_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25870_ _10860_ registers\[47\]\[62\] _11158_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__mux2_1
XFILLER_41_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24821_ _09615_ registers\[54\]\[48\] _10631_ VGND VGND VPWR VPWR _10640_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34999_ clknet_leaf_308_CLK _03113_ VGND VGND VPWR VPWR registers\[21\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27540_ _12137_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__clkbuf_1
X_24752_ _09546_ registers\[54\]\[15\] _10598_ VGND VGND VPWR VPWR _10604_ sky130_fd_sc_hd__mux2_1
X_21964_ registers\[20\]\[36\] registers\[21\]\[36\] registers\[22\]\[36\] registers\[23\]\[36\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__mux4_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23703_ _09510_ registers\[29\]\[0\] _10017_ VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__mux2_1
X_20915_ _07358_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__buf_6
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24683_ _10566_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27471_ _12101_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21895_ _08423_ _08558_ _08559_ _08428_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__a22o_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29210_ net47 VGND VGND VPWR VPWR _13042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26422_ _10737_ registers\[42\]\[3\] _11514_ VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__mux2_1
X_23634_ registers\[61\]\[33\] _09760_ _09976_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__mux2_1
X_20846_ _07536_ _07539_ _07310_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__o21ba_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29141_ net22 VGND VGND VPWR VPWR _12995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_211_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23565_ registers\[61\]\[0\] _09648_ _09943_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__mux2_1
XFILLER_23_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26353_ _11481_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__clkbuf_1
X_20777_ registers\[44\]\[3\] registers\[45\]\[3\] registers\[46\]\[3\] registers\[47\]\[3\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__mux4_1
XFILLER_204_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25304_ _10844_ registers\[51\]\[54\] _10920_ VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__mux2_1
X_22516_ _09012_ _09161_ _09162_ _09018_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__a22o_1
XFILLER_161_1156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26284_ _11445_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29072_ _12948_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__clkbuf_1
X_23496_ _09906_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28023_ _12392_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__clkbuf_1
X_22447_ _07358_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__buf_4
X_25235_ _10775_ registers\[51\]\[21\] _10887_ VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__mux2_1
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25166_ _10848_ registers\[52\]\[56\] _10836_ VGND VGND VPWR VPWR _10849_ sky130_fd_sc_hd__mux2_1
X_22378_ _08953_ _09027_ _09028_ _08956_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__a22o_1
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24117_ _09521_ registers\[58\]\[3\] _10233_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__mux2_1
XFILLER_191_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21329_ registers\[28\]\[18\] registers\[29\]\[18\] registers\[30\]\[18\] registers\[31\]\[18\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__mux4_1
XFILLER_151_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25097_ net28 VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__buf_2
X_29974_ registers\[17\]\[23\] _12983_ _13446_ VGND VGND VPWR VPWR _13450_ sky130_fd_sc_hd__mux2_1
X_28925_ registers\[24\]\[5\] _10315_ _12861_ VGND VGND VPWR VPWR _12867_ sky130_fd_sc_hd__mux2_1
X_24048_ _09588_ registers\[5\]\[35\] _10194_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__mux2_1
XFILLER_133_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16870_ registers\[16\]\[22\] registers\[17\]\[22\] registers\[18\]\[22\] registers\[19\]\[22\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15362_ sky130_fd_sc_hd__mux4_1
X_28856_ _12830_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27807_ registers\[33\]\[51\] _10412_ _12277_ VGND VGND VPWR VPWR _12279_ sky130_fd_sc_hd__mux2_1
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28787_ _12794_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__clkbuf_1
X_25999_ _10854_ registers\[46\]\[59\] _11285_ VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__mux2_1
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18540_ registers\[40\]\[5\] registers\[41\]\[5\] registers\[42\]\[5\] registers\[43\]\[5\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__mux4_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27738_ _12242_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__clkbuf_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _05226_ _05231_ _05163_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__o21ba_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27669_ _12150_ VGND VGND VPWR VPWR _12206_ sky130_fd_sc_hd__buf_4
XFILLER_205_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29408_ _13152_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_352 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17422_ _15891_ _15897_ _15620_ _15621_ VGND VGND VPWR VPWR _15898_ sky130_fd_sc_hd__o211a_1
XANTENNA_363 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30680_ _13821_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_396 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29339_ _09780_ registers\[22\]\[42\] _13113_ VGND VGND VPWR VPWR _13116_ sky130_fd_sc_hd__mux2_1
X_17353_ registers\[12\]\[36\] registers\[13\]\[36\] registers\[14\]\[36\] registers\[15\]\[36\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15831_ sky130_fd_sc_hd__mux4_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16304_ registers\[28\]\[6\] registers\[29\]\[6\] registers\[30\]\[6\] registers\[31\]\[6\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14812_ sky130_fd_sc_hd__mux4_1
X_32350_ clknet_leaf_46_CLK _00464_ VGND VGND VPWR VPWR registers\[61\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17284_ registers\[12\]\[34\] registers\[13\]\[34\] registers\[14\]\[34\] registers\[15\]\[34\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15764_ sky130_fd_sc_hd__mux4_1
XFILLER_173_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19023_ registers\[4\]\[18\] registers\[5\]\[18\] registers\[6\]\[18\] registers\[7\]\[18\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__mux4_1
X_31301_ _14148_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__clkbuf_1
X_16235_ registers\[20\]\[4\] registers\[21\]\[4\] registers\[22\]\[4\] registers\[23\]\[4\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14745_ sky130_fd_sc_hd__mux4_1
XFILLER_139_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32281_ clknet_leaf_6_CLK _00395_ VGND VGND VPWR VPWR registers\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34020_ clknet_leaf_440_CLK _02134_ VGND VGND VPWR VPWR registers\[36\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31232_ registers\[8\]\[43\] net38 _14108_ VGND VGND VPWR VPWR _14112_ sky130_fd_sc_hd__mux2_1
XFILLER_6_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16166_ _14592_ VGND VGND VPWR VPWR _14678_ sky130_fd_sc_hd__buf_6
XFILLER_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31163_ registers\[8\]\[10\] net2 _14075_ VGND VGND VPWR VPWR _14076_ sky130_fd_sc_hd__mux2_1
X_16097_ _14610_ VGND VGND VPWR VPWR _14611_ sky130_fd_sc_hd__buf_4
XFILLER_138_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30114_ _13523_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__clkbuf_1
X_19925_ _05078_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__buf_6
XFILLER_138_1169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35971_ clknet_leaf_232_CLK _04085_ VGND VGND VPWR VPWR registers\[6\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31094_ _14039_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_296_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_296_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30045_ registers\[17\]\[57\] _13054_ _13479_ VGND VGND VPWR VPWR _13487_ sky130_fd_sc_hd__mux2_1
X_19856_ registers\[44\]\[42\] registers\[45\]\[42\] registers\[46\]\[42\] registers\[47\]\[42\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__mux4_1
X_34922_ clknet_leaf_453_CLK _03036_ VGND VGND VPWR VPWR registers\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18807_ _05412_ _05556_ _05557_ _05416_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__a22o_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34853_ clknet_leaf_447_CLK _02967_ VGND VGND VPWR VPWR registers\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_19787_ registers\[52\]\[40\] registers\[53\]\[40\] registers\[54\]\[40\] registers\[55\]\[40\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__mux4_1
X_16999_ _14510_ VGND VGND VPWR VPWR _15487_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33804_ clknet_leaf_171_CLK _01918_ VGND VGND VPWR VPWR registers\[40\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_18738_ registers\[12\]\[10\] registers\[13\]\[10\] registers\[14\]\[10\] registers\[15\]\[10\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__mux4_1
X_34784_ clknet_leaf_9_CLK _02898_ VGND VGND VPWR VPWR registers\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31996_ clknet_leaf_27_CLK _00168_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_1
XFILLER_224_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33735_ clknet_leaf_243_CLK _01849_ VGND VGND VPWR VPWR registers\[41\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_18669_ _05127_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__buf_4
X_30947_ registers\[10\]\[36\] _13010_ _13955_ VGND VGND VPWR VPWR _13962_ sky130_fd_sc_hd__mux2_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20700_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__buf_2
XFILLER_184_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33666_ clknet_leaf_249_CLK _01780_ VGND VGND VPWR VPWR registers\[42\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21680_ registers\[16\]\[28\] registers\[17\]\[28\] registers\[18\]\[28\] registers\[19\]\[28\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__mux4_1
X_30878_ registers\[10\]\[3\] _12941_ _13922_ VGND VGND VPWR VPWR _13926_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35405_ clknet_leaf_133_CLK _03519_ VGND VGND VPWR VPWR registers\[15\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20631_ registers\[60\]\[0\] registers\[61\]\[0\] registers\[62\]\[0\] registers\[63\]\[0\]
+ _07327_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__mux4_1
XFILLER_162_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32617_ clknet_leaf_424_CLK _00731_ VGND VGND VPWR VPWR registers\[58\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33597_ clknet_leaf_274_CLK _01711_ VGND VGND VPWR VPWR registers\[43\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_220_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_220_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35336_ clknet_leaf_154_CLK _03450_ VGND VGND VPWR VPWR registers\[16\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_23350_ registers\[39\]\[29\] _09751_ _09700_ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__mux2_1
X_20562_ registers\[12\]\[63\] registers\[13\]\[63\] registers\[14\]\[63\] registers\[15\]\[63\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__mux4_1
X_32548_ clknet_leaf_470_CLK _00662_ VGND VGND VPWR VPWR registers\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22301_ registers\[8\]\[46\] registers\[9\]\[46\] registers\[10\]\[46\] registers\[11\]\[46\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__mux4_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35267_ clknet_leaf_223_CLK _03381_ VGND VGND VPWR VPWR registers\[17\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_23281_ registers\[9\]\[43\] _09782_ _09776_ VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__mux2_1
X_20493_ registers\[48\]\[61\] registers\[49\]\[61\] registers\[50\]\[61\] registers\[51\]\[61\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__mux4_1
X_32479_ clknet_leaf_48_CLK _00593_ VGND VGND VPWR VPWR registers\[60\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25020_ _10749_ registers\[52\]\[9\] _10731_ VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__mux2_1
XFILLER_146_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22232_ _08677_ _08885_ _08886_ _08681_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__a22o_1
X_34218_ clknet_leaf_427_CLK _02332_ VGND VGND VPWR VPWR registers\[33\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35198_ clknet_leaf_191_CLK _03312_ VGND VGND VPWR VPWR registers\[18\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22163_ _08669_ _08818_ _08819_ _08675_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__a22o_1
X_34149_ clknet_leaf_56_CLK _02263_ VGND VGND VPWR VPWR registers\[34\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21114_ _07586_ _07799_ _07800_ _07589_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__a22o_1
XTAP_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26971_ net43 VGND VGND VPWR VPWR _11830_ sky130_fd_sc_hd__buf_4
X_22094_ _07358_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__buf_4
XTAP_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_287_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_287_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28710_ _11795_ registers\[26\]\[31\] _12752_ VGND VGND VPWR VPWR _12754_ sky130_fd_sc_hd__mux2_1
X_25922_ _10777_ registers\[46\]\[22\] _11252_ VGND VGND VPWR VPWR _11255_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21045_ registers\[16\]\[10\] registers\[17\]\[10\] registers\[18\]\[10\] registers\[19\]\[10\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__mux4_1
X_29690_ _13300_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28641_ _11861_ registers\[27\]\[63\] _12647_ VGND VGND VPWR VPWR _12717_ sky130_fd_sc_hd__mux2_1
X_25853_ _11218_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24804_ _10586_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__buf_4
XFILLER_46_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28572_ _12647_ VGND VGND VPWR VPWR _12681_ sky130_fd_sc_hd__buf_4
XFILLER_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25784_ _11182_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22996_ _09593_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27523_ _12128_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24735_ _09529_ registers\[54\]\[7\] _10587_ VGND VGND VPWR VPWR _10595_ sky130_fd_sc_hd__mux2_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21947_ _07275_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__buf_4
XFILLER_216_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27454_ _12092_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21878_ registers\[52\]\[34\] registers\[53\]\[34\] registers\[54\]\[34\] registers\[55\]\[34\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__mux4_1
X_24666_ _10557_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26405_ _11508_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__clkbuf_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20829_ _07347_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__buf_6
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ registers\[61\]\[25\] _09742_ _09965_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__mux2_1
XFILLER_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27385_ registers\[36\]\[44\] _10397_ _12051_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__mux2_1
X_24597_ _10521_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_211_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_211_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_29124_ registers\[23\]\[23\] _12983_ _12977_ VGND VGND VPWR VPWR _12984_ sky130_fd_sc_hd__mux2_1
X_26336_ _11472_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23548_ _09933_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29055_ net12 VGND VGND VPWR VPWR _12937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26267_ _10852_ registers\[44\]\[58\] _11427_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__mux2_1
X_23479_ _09897_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16020_ _14493_ VGND VGND VPWR VPWR _14534_ sky130_fd_sc_hd__buf_4
X_28006_ _12383_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25218_ _10758_ registers\[51\]\[13\] _10876_ VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26198_ _10783_ registers\[44\]\[25\] _11394_ VGND VGND VPWR VPWR _11400_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25149_ _10837_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17971_ registers\[40\]\[54\] registers\[41\]\[54\] registers\[42\]\[54\] registers\[43\]\[54\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux4_1
XFILLER_3_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29957_ registers\[17\]\[15\] _12966_ _13435_ VGND VGND VPWR VPWR _13441_ sky130_fd_sc_hd__mux2_1
XFILLER_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_278_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_278_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19710_ registers\[56\]\[38\] registers\[57\]\[38\] registers\[58\]\[38\] registers\[59\]\[38\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__mux4_1
X_28908_ _12857_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__clkbuf_1
X_16922_ _15198_ _15410_ _15411_ _15204_ VGND VGND VPWR VPWR _15412_ sky130_fd_sc_hd__a22o_1
X_29888_ _13404_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19641_ registers\[60\]\[36\] registers\[61\]\[36\] registers\[62\]\[36\] registers\[63\]\[36\]
+ _06305_ _06099_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__mux4_1
XFILLER_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28839_ _12821_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16853_ _15341_ _15342_ _15343_ _15344_ VGND VGND VPWR VPWR _15345_ sky130_fd_sc_hd__a22o_1
XFILLER_172_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19572_ _05078_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__buf_6
X_31850_ _09691_ registers\[49\]\[16\] _14430_ VGND VGND VPWR VPWR _14437_ sky130_fd_sc_hd__mux2_1
X_16784_ _14555_ VGND VGND VPWR VPWR _15278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_219_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18523_ registers\[0\]\[4\] registers\[1\]\[4\] registers\[2\]\[4\] registers\[3\]\[4\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__mux4_1
X_30801_ _13885_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31781_ _14400_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33520_ clknet_leaf_361_CLK _01634_ VGND VGND VPWR VPWR registers\[44\]\[34\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_450_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_450_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30732_ _13848_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__clkbuf_1
X_18454_ _05089_ _05213_ _05214_ _05100_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a22o_1
XFILLER_146_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_182 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ registers\[36\]\[38\] registers\[37\]\[38\] registers\[38\]\[38\] registers\[39\]\[38\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _15881_ sky130_fd_sc_hd__mux4_1
XANTENNA_193 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33451_ clknet_leaf_429_CLK _01565_ VGND VGND VPWR VPWR registers\[45\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18385_ _05137_ _05140_ _05145_ _05147_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__a22o_1
XFILLER_18_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30663_ _13812_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__clkbuf_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_202_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_202_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32402_ clknet_leaf_101_CLK _00516_ VGND VGND VPWR VPWR registers\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36170_ clknet_leaf_177_CLK _04284_ VGND VGND VPWR VPWR registers\[49\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_17336_ _15684_ _15812_ _15813_ _15687_ VGND VGND VPWR VPWR _15814_ sky130_fd_sc_hd__a22o_1
XFILLER_159_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33382_ clknet_leaf_58_CLK _01496_ VGND VGND VPWR VPWR registers\[46\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_30594_ _09821_ registers\[13\]\[61\] _13708_ VGND VGND VPWR VPWR _13776_ sky130_fd_sc_hd__mux2_1
XFILLER_202_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35121_ clknet_leaf_381_CLK _03235_ VGND VGND VPWR VPWR registers\[1\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_32333_ clknet_leaf_144_CLK _00447_ VGND VGND VPWR VPWR registers\[19\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17267_ _15677_ _15745_ _15746_ _15682_ VGND VGND VPWR VPWR _15747_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19006_ _05045_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__clkbuf_4
X_16218_ registers\[60\]\[4\] registers\[61\]\[4\] registers\[62\]\[4\] registers\[63\]\[4\]
+ _14727_ _14544_ VGND VGND VPWR VPWR _14728_ sky130_fd_sc_hd__mux4_1
XFILLER_128_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35052_ clknet_leaf_395_CLK _03166_ VGND VGND VPWR VPWR registers\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_32264_ clknet_leaf_237_CLK _00378_ VGND VGND VPWR VPWR registers\[39\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17198_ registers\[40\]\[32\] registers\[41\]\[32\] registers\[42\]\[32\] registers\[43\]\[32\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15680_ sky130_fd_sc_hd__mux4_1
X_34003_ clknet_leaf_127_CLK _02117_ VGND VGND VPWR VPWR registers\[36\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_31215_ registers\[8\]\[35\] net29 _14097_ VGND VGND VPWR VPWR _14103_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16149_ registers\[56\]\[2\] registers\[57\]\[2\] registers\[58\]\[2\] registers\[59\]\[2\]
+ _14530_ _14532_ VGND VGND VPWR VPWR _14661_ sky130_fd_sc_hd__mux4_1
XFILLER_161_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32195_ clknet_leaf_399_CLK _00309_ VGND VGND VPWR VPWR registers\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31146_ registers\[8\]\[2\] net23 _14064_ VGND VGND VPWR VPWR _14067_ sky130_fd_sc_hd__mux2_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_269_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_269_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_233_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19908_ _06622_ _06627_ _06523_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__o21ba_1
XFILLER_229_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31077_ _14030_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__clkbuf_1
X_35954_ clknet_leaf_380_CLK _04068_ VGND VGND VPWR VPWR registers\[6\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30028_ registers\[17\]\[49\] _13037_ _13468_ VGND VGND VPWR VPWR _13478_ sky130_fd_sc_hd__mux2_1
X_34905_ clknet_leaf_4_CLK _03019_ VGND VGND VPWR VPWR registers\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19839_ registers\[24\]\[41\] registers\[25\]\[41\] registers\[26\]\[41\] registers\[27\]\[41\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__mux4_1
XFILLER_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35885_ clknet_leaf_391_CLK _03999_ VGND VGND VPWR VPWR registers\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22850_ _07325_ _09484_ _09485_ _07336_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__a22o_1
X_34836_ clknet_leaf_98_CLK _02950_ VGND VGND VPWR VPWR registers\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21801_ _08462_ _08465_ _08466_ _08467_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__a22o_1
X_22781_ _07355_ _09418_ _09419_ _07367_ VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__a22o_1
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34767_ clknet_leaf_111_CLK _02881_ VGND VGND VPWR VPWR registers\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_31979_ clknet_leaf_21_CLK _00149_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_224_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_441_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_441_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24520_ _10479_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
X_21732_ _08326_ _08399_ _08400_ _08332_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__a22o_1
X_33718_ clknet_leaf_341_CLK _01832_ VGND VGND VPWR VPWR registers\[41\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_34698_ clknet_leaf_152_CLK _02812_ VGND VGND VPWR VPWR registers\[26\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24451_ _10443_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
X_21663_ _07324_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__clkbuf_8
XFILLER_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33649_ clknet_leaf_347_CLK _01763_ VGND VGND VPWR VPWR registers\[42\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23402_ _09855_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
X_20614_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27170_ _11742_ registers\[37\]\[6\] _11936_ VGND VGND VPWR VPWR _11943_ sky130_fd_sc_hd__mux2_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24382_ net39 VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21594_ _07275_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__buf_4
XFILLER_36_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23333_ net55 VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__buf_4
X_26121_ _11359_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
X_20545_ registers\[40\]\[63\] registers\[41\]\[63\] registers\[42\]\[63\] registers\[43\]\[63\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__mux4_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35319_ clknet_leaf_311_CLK _03433_ VGND VGND VPWR VPWR registers\[16\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26052_ _11300_ VGND VGND VPWR VPWR _11323_ sky130_fd_sc_hd__buf_4
X_23264_ net32 VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__clkbuf_4
X_20476_ registers\[24\]\[60\] registers\[25\]\[60\] registers\[26\]\[60\] registers\[27\]\[60\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__mux4_1
XFILLER_180_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25003_ _10738_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
X_22215_ _08867_ _08870_ _08773_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__o21ba_1
X_23195_ registers\[9\]\[15\] _09689_ _09722_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29811_ _13352_ VGND VGND VPWR VPWR _13364_ sky130_fd_sc_hd__buf_4
XTAP_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22146_ _08782_ _08789_ _08796_ _08803_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__or4_4
XTAP_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1509 _07395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29742_ registers\[1\]\[41\] _13021_ _13326_ VGND VGND VPWR VPWR _13328_ sky130_fd_sc_hd__mux2_1
XTAP_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26954_ _11818_ registers\[3\]\[42\] _11814_ VGND VGND VPWR VPWR _11819_ sky130_fd_sc_hd__mux2_1
X_22077_ _07333_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__clkbuf_4
XTAP_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21028_ registers\[52\]\[10\] registers\[53\]\[10\] registers\[54\]\[10\] registers\[55\]\[10\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__mux4_1
X_25905_ _10760_ registers\[46\]\[14\] _11241_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__mux2_1
X_29673_ _13291_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26885_ _11729_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__buf_4
XFILLER_43_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28624_ _12708_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__clkbuf_1
X_25836_ _11209_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28555_ _12672_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25767_ _11173_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22979_ net26 VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__clkbuf_4
XFILLER_231_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_432_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_432_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27506_ _12119_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__clkbuf_1
X_24718_ _09511_ _10584_ VGND VGND VPWR VPWR _10585_ sky130_fd_sc_hd__nor2_8
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28486_ _11841_ registers\[28\]\[53\] _12632_ VGND VGND VPWR VPWR _12636_ sky130_fd_sc_hd__mux2_1
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25698_ registers\[48\]\[45\] _10399_ _11130_ VGND VGND VPWR VPWR _11136_ sky130_fd_sc_hd__mux2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27437_ _12083_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__clkbuf_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _09580_ registers\[55\]\[31\] _10547_ VGND VGND VPWR VPWR _10549_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ registers\[0\]\[60\] registers\[1\]\[60\] registers\[2\]\[60\] registers\[3\]\[60\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__mux4_1
X_27368_ registers\[36\]\[36\] _10380_ _12040_ VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29107_ net10 VGND VGND VPWR VPWR _12972_ sky130_fd_sc_hd__clkbuf_4
X_17121_ registers\[32\]\[30\] registers\[33\]\[30\] registers\[34\]\[30\] registers\[35\]\[30\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15605_ sky130_fd_sc_hd__mux4_1
X_26319_ _11463_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
X_27299_ registers\[36\]\[3\] _10311_ _12007_ VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__mux2_1
XFILLER_7_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_35__f_CLK clknet_5_17_0_CLK VGND VGND VPWR VPWR clknet_6_35__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29038_ registers\[24\]\[59\] _10428_ _12916_ VGND VGND VPWR VPWR _12926_ sky130_fd_sc_hd__mux2_1
XFILLER_128_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17052_ registers\[36\]\[28\] registers\[37\]\[28\] registers\[38\]\[28\] registers\[39\]\[28\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15538_ sky130_fd_sc_hd__mux4_1
XFILLER_183_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16003_ _14516_ VGND VGND VPWR VPWR _14517_ sky130_fd_sc_hd__buf_4
XFILLER_100_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31000_ _13989_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17954_ registers\[0\]\[53\] registers\[1\]\[53\] registers\[2\]\[53\] registers\[3\]\[53\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__mux4_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16905_ _15290_ _15394_ _15395_ _15293_ VGND VGND VPWR VPWR _15396_ sky130_fd_sc_hd__a22o_1
XFILLER_61_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32951_ clknet_leaf_327_CLK _01065_ VGND VGND VPWR VPWR registers\[53\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_17885_ registers\[8\]\[51\] registers\[9\]\[51\] registers\[10\]\[51\] registers\[11\]\[51\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31902_ _14464_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19624_ _06182_ _06350_ _06351_ _06185_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__a22o_1
X_16836_ registers\[28\]\[21\] registers\[29\]\[21\] registers\[30\]\[21\] registers\[31\]\[21\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15329_ sky130_fd_sc_hd__mux4_1
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35670_ clknet_leaf_86_CLK _03784_ VGND VGND VPWR VPWR registers\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_32882_ clknet_leaf_356_CLK _00996_ VGND VGND VPWR VPWR registers\[54\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34621_ clknet_leaf_182_CLK _02735_ VGND VGND VPWR VPWR registers\[27\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31833_ _09674_ registers\[49\]\[8\] _14419_ VGND VGND VPWR VPWR _14428_ sky130_fd_sc_hd__mux2_1
X_19555_ _06279_ _06284_ _06180_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__o21ba_1
XFILLER_207_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16767_ registers\[40\]\[20\] registers\[41\]\[20\] registers\[42\]\[20\] registers\[43\]\[20\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15261_ sky130_fd_sc_hd__mux4_1
XFILLER_202_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18506_ registers\[40\]\[4\] registers\[41\]\[4\] registers\[42\]\[4\] registers\[43\]\[4\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__mux4_1
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_423_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_423_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_207_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34552_ clknet_leaf_309_CLK _02666_ VGND VGND VPWR VPWR registers\[28\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19486_ registers\[24\]\[31\] registers\[25\]\[31\] registers\[26\]\[31\] registers\[27\]\[31\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__mux4_1
X_31764_ _14391_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__clkbuf_1
X_16698_ registers\[44\]\[18\] registers\[45\]\[18\] registers\[46\]\[18\] registers\[47\]\[18\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15194_ sky130_fd_sc_hd__mux4_1
XFILLER_206_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30715_ registers\[12\]\[54\] _13048_ _13835_ VGND VGND VPWR VPWR _13840_ sky130_fd_sc_hd__mux2_1
XFILLER_179_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18437_ _05042_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__buf_6
XFILLER_59_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33503_ clknet_leaf_39_CLK _01617_ VGND VGND VPWR VPWR registers\[44\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_34483_ clknet_leaf_384_CLK _02597_ VGND VGND VPWR VPWR registers\[2\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31695_ _14355_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__clkbuf_1
X_36222_ clknet_leaf_116_CLK _00106_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dfxtp_1
X_33434_ clknet_leaf_31_CLK _01548_ VGND VGND VPWR VPWR registers\[45\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_18368_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__clkbuf_4
X_30646_ registers\[12\]\[21\] _12979_ _13802_ VGND VGND VPWR VPWR _13804_ sky130_fd_sc_hd__mux2_1
X_36153_ clknet_leaf_281_CLK _04267_ VGND VGND VPWR VPWR registers\[49\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17319_ registers\[4\]\[35\] registers\[5\]\[35\] registers\[6\]\[35\] registers\[7\]\[35\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15798_ sky130_fd_sc_hd__mux4_1
X_33365_ clknet_leaf_123_CLK _01479_ VGND VGND VPWR VPWR registers\[46\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18299_ _05053_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__clkbuf_4
X_30577_ _13767_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20330_ registers\[20\]\[55\] registers\[21\]\[55\] registers\[22\]\[55\] registers\[23\]\[55\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__mux4_1
X_32316_ clknet_leaf_190_CLK _00430_ VGND VGND VPWR VPWR registers\[19\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_35104_ clknet_leaf_485_CLK _03218_ VGND VGND VPWR VPWR registers\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_36084_ clknet_leaf_351_CLK _04198_ VGND VGND VPWR VPWR registers\[59\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_33296_ clknet_leaf_129_CLK _01410_ VGND VGND VPWR VPWR registers\[47\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35035_ clknet_leaf_492_CLK _03149_ VGND VGND VPWR VPWR registers\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20261_ _06965_ _06970_ _06866_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__o21ba_1
X_32247_ clknet_leaf_336_CLK _00361_ VGND VGND VPWR VPWR registers\[39\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22000_ _08661_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__buf_6
XFILLER_66_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20192_ registers\[24\]\[51\] registers\[25\]\[51\] registers\[26\]\[51\] registers\[27\]\[51\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__mux4_1
XFILLER_118_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32178_ clknet_leaf_14_CLK _00292_ VGND VGND VPWR VPWR registers\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31129_ _14057_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__clkbuf_1
XTAP_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _10148_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35937_ clknet_leaf_481_CLK _04051_ VGND VGND VPWR VPWR registers\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22902_ _09529_ registers\[62\]\[7\] _09515_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__mux2_1
X_26670_ _11648_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35868_ clknet_leaf_478_CLK _03982_ VGND VGND VPWR VPWR registers\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_23882_ _10112_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
X_25621_ _11095_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
X_34819_ clknet_leaf_224_CLK _02933_ VGND VGND VPWR VPWR registers\[24\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_22833_ registers\[4\]\[62\] registers\[5\]\[62\] registers\[6\]\[62\] registers\[7\]\[62\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__mux4_1
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_907 _09681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_918 _09758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35799_ clknet_leaf_85_CLK _03913_ VGND VGND VPWR VPWR registers\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_929 _09869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_414_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_414_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28340_ registers\[2\]\[48\] _10405_ _12550_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25552_ registers\[4\]\[41\] _10391_ _11056_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__mux2_1
X_22764_ _07372_ _09401_ _09402_ _07382_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__a22o_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24503_ _10470_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21715_ registers\[20\]\[29\] registers\[21\]\[29\] registers\[22\]\[29\] registers\[23\]\[29\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__mux4_1
X_28271_ registers\[2\]\[15\] _10336_ _12517_ VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22695_ registers\[40\]\[58\] registers\[41\]\[58\] registers\[42\]\[58\] registers\[43\]\[58\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__mux4_1
X_25483_ _11021_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27222_ _11970_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__clkbuf_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24434_ net58 VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_205_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21646_ _08296_ _08303_ _08310_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__or4_4
XFILLER_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27153_ _11933_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__clkbuf_1
X_21577_ _08250_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
X_24365_ _10385_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_60 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26104_ _11350_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_82 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23316_ net50 VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__buf_4
XANTENNA_93 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20528_ _07225_ _07228_ _05102_ _05104_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__o211a_1
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27084_ _11897_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_1
X_24296_ registers\[57\]\[16\] _10338_ _10326_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__mux2_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26035_ _11314_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20459_ registers\[36\]\[60\] registers\[37\]\[60\] registers\[38\]\[60\] registers\[39\]\[60\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__mux4_1
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23247_ net27 VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23178_ registers\[9\]\[7\] _09672_ _09709_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__mux2_1
XFILLER_79_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1306 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1317 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22129_ registers\[52\]\[41\] registers\[53\]\[41\] registers\[54\]\[41\] registers\[55\]\[41\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__mux4_1
XTAP_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1328 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27986_ _11746_ registers\[31\]\[8\] _12364_ VGND VGND VPWR VPWR _12373_ sky130_fd_sc_hd__mux2_1
XANTENNA_1339 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29725_ registers\[1\]\[33\] _13004_ _13315_ VGND VGND VPWR VPWR _13319_ sky130_fd_sc_hd__mux2_1
XTAP_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26937_ net31 VGND VGND VPWR VPWR _11807_ sky130_fd_sc_hd__clkbuf_4
XTAP_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29656_ registers\[1\]\[0\] _12931_ _13282_ VGND VGND VPWR VPWR _13283_ sky130_fd_sc_hd__mux2_1
X_17670_ _15825_ _04450_ _04451_ _15828_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__a22o_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26868_ _11760_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28607_ _12699_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__clkbuf_1
X_16621_ _14952_ _15118_ _15119_ _14957_ VGND VGND VPWR VPWR _15120_ sky130_fd_sc_hd__a22o_1
XFILLER_60_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25819_ _11200_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
X_29587_ _13246_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__clkbuf_1
X_26799_ registers\[40\]\[53\] _10416_ _11713_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_405_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_405_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19340_ registers\[16\]\[27\] registers\[17\]\[27\] registers\[18\]\[27\] registers\[19\]\[27\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__mux4_1
XFILLER_1_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16552_ _14947_ _15051_ _15052_ _14950_ VGND VGND VPWR VPWR _15053_ sky130_fd_sc_hd__a22o_1
X_28538_ _12663_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19271_ _05839_ _06007_ _06008_ _05842_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a22o_1
X_28469_ _11824_ registers\[28\]\[45\] _12621_ VGND VGND VPWR VPWR _12627_ sky130_fd_sc_hd__mux2_1
X_16483_ registers\[28\]\[11\] registers\[29\]\[11\] registers\[30\]\[11\] registers\[31\]\[11\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14986_ sky130_fd_sc_hd__mux4_1
XFILLER_203_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18222_ registers\[56\]\[62\] registers\[57\]\[62\] registers\[58\]\[62\] registers\[59\]\[62\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__mux4_1
X_30500_ _09691_ registers\[13\]\[16\] _13720_ VGND VGND VPWR VPWR _13727_ sky130_fd_sc_hd__mux2_1
XFILLER_231_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31480_ _14242_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18153_ _04899_ _04906_ _04913_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__or4_4
X_30431_ _13690_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17104_ registers\[8\]\[29\] registers\[9\]\[29\] registers\[10\]\[29\] registers\[11\]\[29\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15589_ sky130_fd_sc_hd__mux4_1
X_33150_ clknet_leaf_268_CLK _01264_ VGND VGND VPWR VPWR registers\[50\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_18084_ _14511_ _04852_ _04853_ _14517_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__a22o_1
X_30362_ _13654_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32101_ clknet_leaf_483_CLK _00015_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dfxtp_1
XFILLER_144_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17035_ registers\[12\]\[27\] registers\[13\]\[27\] registers\[14\]\[27\] registers\[15\]\[27\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15522_ sky130_fd_sc_hd__mux4_1
X_33081_ clknet_leaf_285_CLK _01195_ VGND VGND VPWR VPWR registers\[51\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_30293_ _13617_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32032_ clknet_leaf_44_CLK _00210_ VGND VGND VPWR VPWR registers\[62\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ registers\[24\]\[17\] registers\[25\]\[17\] registers\[26\]\[17\] registers\[27\]\[17\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__mux4_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17937_ _04688_ _04695_ _04702_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__or4_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33983_ clknet_leaf_269_CLK _02097_ VGND VGND VPWR VPWR registers\[37\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35722_ clknet_leaf_153_CLK _03836_ VGND VGND VPWR VPWR registers\[10\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17868_ _04636_ _04643_ _04644_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__o21ba_1
X_32934_ clknet_leaf_437_CLK _01048_ VGND VGND VPWR VPWR registers\[53\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19607_ registers\[48\]\[35\] registers\[49\]\[35\] registers\[50\]\[35\] registers\[51\]\[35\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__mux4_1
X_35653_ clknet_leaf_214_CLK _03767_ VGND VGND VPWR VPWR registers\[11\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_16819_ registers\[56\]\[21\] registers\[57\]\[21\] registers\[58\]\[21\] registers\[59\]\[21\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15312_ sky130_fd_sc_hd__mux4_1
XFILLER_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17799_ registers\[44\]\[49\] registers\[45\]\[49\] registers\[46\]\[49\] registers\[47\]\[49\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__mux4_1
X_32865_ clknet_leaf_44_CLK _00979_ VGND VGND VPWR VPWR registers\[54\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34604_ clknet_leaf_410_CLK _02718_ VGND VGND VPWR VPWR registers\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31816_ _14418_ VGND VGND VPWR VPWR _14419_ sky130_fd_sc_hd__buf_4
X_19538_ _06233_ _06266_ _06267_ _06236_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__a22o_1
X_35584_ clknet_leaf_237_CLK _03698_ VGND VGND VPWR VPWR registers\[12\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_32796_ clknet_leaf_52_CLK _00910_ VGND VGND VPWR VPWR registers\[55\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31747_ registers\[59\]\[31\] net25 _14381_ VGND VGND VPWR VPWR _14383_ sky130_fd_sc_hd__mux2_1
X_34535_ clknet_leaf_456_CLK _02649_ VGND VGND VPWR VPWR registers\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_19469_ registers\[36\]\[31\] registers\[37\]\[31\] registers\[38\]\[31\] registers\[39\]\[31\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__mux4_1
X_21500_ registers\[4\]\[23\] registers\[5\]\[23\] registers\[6\]\[23\] registers\[7\]\[23\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__mux4_1
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22480_ _09012_ _09126_ _09127_ _09018_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__a22o_1
X_31678_ registers\[63\]\[63\] net60 _14276_ VGND VGND VPWR VPWR _14346_ sky130_fd_sc_hd__mux2_1
X_34466_ clknet_leaf_466_CLK _02580_ VGND VGND VPWR VPWR registers\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36205_ clknet_leaf_100_CLK _00088_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dfxtp_1
X_21431_ _07929_ _08107_ _08108_ _07932_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__a22o_1
X_33417_ clknet_leaf_254_CLK _01531_ VGND VGND VPWR VPWR registers\[46\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_30629_ registers\[12\]\[13\] _12962_ _13791_ VGND VGND VPWR VPWR _13795_ sky130_fd_sc_hd__mux2_1
XFILLER_198_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34397_ clknet_leaf_492_CLK _02511_ VGND VGND VPWR VPWR registers\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24150_ _09554_ registers\[58\]\[19\] _10244_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__mux2_1
X_33348_ clknet_leaf_251_CLK _01462_ VGND VGND VPWR VPWR registers\[47\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_21362_ registers\[20\]\[19\] registers\[21\]\[19\] registers\[22\]\[19\] registers\[23\]\[19\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__mux4_1
X_36136_ clknet_leaf_435_CLK _04250_ VGND VGND VPWR VPWR registers\[49\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23101_ _09667_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
X_20313_ registers\[48\]\[55\] registers\[49\]\[55\] registers\[50\]\[55\] registers\[51\]\[55\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__mux4_1
XFILLER_107_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24081_ _10217_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
Xinput80 R3[3] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
X_33279_ clknet_leaf_268_CLK _01393_ VGND VGND VPWR VPWR registers\[48\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_36067_ clknet_leaf_443_CLK _04181_ VGND VGND VPWR VPWR registers\[59\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_21293_ _07953_ _07960_ _07967_ _07974_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__or4_2
X_23032_ _09617_ registers\[62\]\[49\] _09599_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__mux2_1
X_35018_ clknet_leaf_142_CLK _03132_ VGND VGND VPWR VPWR registers\[21\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_20244_ _06919_ _06952_ _06953_ _06922_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__a22o_1
XFILLER_66_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27840_ _12296_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__clkbuf_1
X_20175_ registers\[36\]\[51\] registers\[37\]\[51\] registers\[38\]\[51\] registers\[39\]\[51\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__mux4_1
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27771_ registers\[33\]\[34\] _10376_ _12255_ VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__mux2_1
X_24983_ _09642_ registers\[53\]\[61\] _10657_ VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__mux2_1
XFILLER_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29510_ _13205_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__clkbuf_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26722_ _11676_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_1
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _10139_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29441_ _13169_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__clkbuf_1
X_26653_ _11639_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_1
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_704 _07285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23865_ _10103_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_715 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25604_ registers\[48\]\[0\] _10303_ _11086_ VGND VGND VPWR VPWR _11087_ sky130_fd_sc_hd__mux2_1
XANTENNA_726 _07349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29372_ _09815_ registers\[22\]\[58\] _13124_ VGND VGND VPWR VPWR _13133_ sky130_fd_sc_hd__mux2_1
X_22816_ registers\[32\]\[62\] registers\[33\]\[62\] registers\[34\]\[62\] registers\[35\]\[62\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__mux4_1
XANTENNA_737 _07358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26584_ _11603_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_748 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23796_ _10066_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_759 _07398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28323_ _12505_ VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__buf_4
XFILLER_246_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25535_ registers\[4\]\[33\] _10374_ _11045_ VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__mux2_1
X_22747_ registers\[16\]\[59\] registers\[17\]\[59\] registers\[18\]\[59\] registers\[19\]\[59\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__mux4_1
XFILLER_198_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28254_ registers\[2\]\[7\] _10319_ _12506_ VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__mux2_1
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25466_ registers\[4\]\[0\] _10303_ _11012_ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__mux2_1
XFILLER_158_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22678_ _09316_ _09319_ _09091_ _09092_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__o211a_1
XFILLER_200_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27205_ _11961_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__clkbuf_1
X_24417_ registers\[57\]\[55\] _10420_ _10410_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21629_ registers\[52\]\[27\] registers\[53\]\[27\] registers\[54\]\[27\] registers\[55\]\[27\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__mux4_1
X_28185_ _12477_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25397_ _10974_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27136_ _11843_ registers\[38\]\[54\] _11920_ VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24348_ net27 VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__buf_4
XFILLER_10_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27067_ _11774_ registers\[38\]\[21\] _11887_ VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__mux2_1
X_24279_ _10327_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_21_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_21_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26018_ _11305_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1103 _14546_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1114 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18840_ _05586_ _05589_ _05483_ _05484_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__o211a_2
XFILLER_49_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1125 _14584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1136 _14613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1147 _15572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18771_ _05412_ _05521_ _05522_ _05416_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1158 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27969_ _12363_ VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__buf_4
X_15983_ _14496_ VGND VGND VPWR VPWR _14497_ sky130_fd_sc_hd__clkbuf_8
XTAP_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1169 _15744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ registers\[40\]\[47\] registers\[41\]\[47\] registers\[42\]\[47\] registers\[43\]\[47\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__mux4_1
XTAP_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29708_ registers\[1\]\[25\] _12987_ _13304_ VGND VGND VPWR VPWR _13310_ sky130_fd_sc_hd__mux2_1
X_30980_ _13979_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__clkbuf_1
XTAP_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ registers\[32\]\[45\] registers\[33\]\[45\] registers\[34\]\[45\] registers\[35\]\[45\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__mux4_1
XFILLER_110_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29639_ _13273_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__clkbuf_1
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16604_ registers\[52\]\[15\] registers\[53\]\[15\] registers\[54\]\[15\] registers\[55\]\[15\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _15103_ sky130_fd_sc_hd__mux4_1
X_32650_ clknet_leaf_176_CLK _00764_ VGND VGND VPWR VPWR registers\[58\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17584_ _04345_ _04352_ _04359_ _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__or4_1
XFILLER_21_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31601_ registers\[63\]\[26\] net19 _14299_ VGND VGND VPWR VPWR _14306_ sky130_fd_sc_hd__mux2_1
X_19323_ _05890_ _06055_ _06058_ _05893_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__a22o_1
XFILLER_91_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16535_ registers\[48\]\[13\] registers\[49\]\[13\] registers\[50\]\[13\] registers\[51\]\[13\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15036_ sky130_fd_sc_hd__mux4_1
X_32581_ clknet_leaf_232_CLK _00695_ VGND VGND VPWR VPWR registers\[5\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31532_ _14269_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__clkbuf_1
X_34320_ clknet_leaf_100_CLK _02434_ VGND VGND VPWR VPWR registers\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_19254_ registers\[48\]\[25\] registers\[49\]\[25\] registers\[50\]\[25\] registers\[51\]\[25\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__mux4_1
X_16466_ registers\[56\]\[11\] registers\[57\]\[11\] registers\[58\]\[11\] registers\[59\]\[11\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _14969_ sky130_fd_sc_hd__mux4_1
XFILLER_231_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18205_ _04967_ _04970_ _14584_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__o21ba_1
X_34251_ clknet_leaf_157_CLK _02365_ VGND VGND VPWR VPWR registers\[33\]\[61\] sky130_fd_sc_hd__dfxtp_1
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31463_ _14233_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__clkbuf_1
X_19185_ _05890_ _05923_ _05924_ _05893_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__a22o_1
X_16397_ _14898_ _14901_ _14554_ _14556_ VGND VGND VPWR VPWR _14902_ sky130_fd_sc_hd__o211a_1
X_33202_ clknet_leaf_379_CLK _01316_ VGND VGND VPWR VPWR registers\[4\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_18136_ registers\[52\]\[59\] registers\[53\]\[59\] registers\[54\]\[59\] registers\[55\]\[59\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux4_1
XFILLER_163_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30414_ _13681_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34182_ clknet_leaf_247_CLK _02296_ VGND VGND VPWR VPWR registers\[34\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31394_ registers\[7\]\[56\] net52 _14190_ VGND VGND VPWR VPWR _14197_ sky130_fd_sc_hd__mux2_1
XFILLER_157_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33133_ clknet_leaf_379_CLK _01247_ VGND VGND VPWR VPWR registers\[50\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_18067_ _04676_ _04835_ _04836_ _04681_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__a22o_1
XFILLER_156_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30345_ _13645_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17018_ _15334_ _15503_ _15504_ _15339_ VGND VGND VPWR VPWR _15505_ sky130_fd_sc_hd__a22o_1
X_33064_ clknet_leaf_435_CLK _01178_ VGND VGND VPWR VPWR registers\[51\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30276_ _13608_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32015_ clknet_leaf_172_CLK _00193_ VGND VGND VPWR VPWR registers\[62\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_916 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18969_ registers\[36\]\[17\] registers\[37\]\[17\] registers\[38\]\[17\] registers\[39\]\[17\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__mux4_1
XFILLER_100_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1670 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1681 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1692 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21980_ _08326_ _08640_ _08641_ _08332_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__a22o_1
X_33966_ clknet_leaf_356_CLK _02080_ VGND VGND VPWR VPWR registers\[37\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35705_ clknet_leaf_317_CLK _03819_ VGND VGND VPWR VPWR registers\[10\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20931_ _07586_ _07621_ _07622_ _07589_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__a22o_1
X_32917_ clknet_leaf_183_CLK _01031_ VGND VGND VPWR VPWR registers\[53\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33897_ clknet_leaf_424_CLK _02011_ VGND VGND VPWR VPWR registers\[38\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20862_ _07552_ _07555_ _07370_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__o21ba_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35636_ clknet_leaf_415_CLK _03750_ VGND VGND VPWR VPWR registers\[11\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_23650_ _09988_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32848_ clknet_leaf_175_CLK _00962_ VGND VGND VPWR VPWR registers\[54\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22601_ _09109_ _09244_ _09245_ _09114_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__a22o_1
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20793_ registers\[12\]\[3\] registers\[13\]\[3\] registers\[14\]\[3\] registers\[15\]\[3\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__mux4_1
X_23581_ registers\[61\]\[8\] _09674_ _09943_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__mux2_1
X_35567_ clknet_leaf_376_CLK _03681_ VGND VGND VPWR VPWR registers\[12\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32779_ clknet_leaf_164_CLK _00893_ VGND VGND VPWR VPWR registers\[56\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25320_ _10860_ registers\[51\]\[62\] _10864_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__mux2_1
XFILLER_50_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22532_ _07363_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__buf_4
X_34518_ clknet_leaf_94_CLK _02632_ VGND VGND VPWR VPWR registers\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35498_ clknet_leaf_398_CLK _03612_ VGND VGND VPWR VPWR registers\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_25251_ _10791_ registers\[51\]\[29\] _10887_ VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__mux2_1
X_34449_ clknet_leaf_106_CLK _02563_ VGND VGND VPWR VPWR registers\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_22463_ _07329_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__buf_4
X_24202_ _10281_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21414_ _07776_ _08090_ _08091_ _07781_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__a22o_1
X_25182_ _10859_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__clkbuf_1
X_22394_ registers\[40\]\[49\] registers\[41\]\[49\] registers\[42\]\[49\] registers\[43\]\[49\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__mux4_1
XFILLER_176_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36119_ clknet_leaf_68_CLK _04233_ VGND VGND VPWR VPWR registers\[49\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_24133_ _10245_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__clkbuf_1
X_21345_ registers\[48\]\[19\] registers\[49\]\[19\] registers\[50\]\[19\] registers\[51\]\[19\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__mux4_1
XFILLER_204_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29990_ _13458_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24064_ _10208_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__clkbuf_1
X_28941_ _12875_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21276_ registers\[52\]\[17\] registers\[53\]\[17\] registers\[54\]\[17\] registers\[55\]\[17\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__mux4_1
XFILLER_144_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20227_ _06934_ _06937_ _06866_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__o21ba_1
X_23015_ _09606_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28872_ _11822_ registers\[25\]\[44\] _12834_ VGND VGND VPWR VPWR _12839_ sky130_fd_sc_hd__mux2_1
XFILLER_85_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27823_ registers\[33\]\[59\] _10428_ _12277_ VGND VGND VPWR VPWR _12287_ sky130_fd_sc_hd__mux2_1
XFILLER_134_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20158_ _05116_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27754_ registers\[33\]\[26\] _10359_ _12244_ VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__mux2_1
XFILLER_218_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24966_ _10716_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__clkbuf_1
X_20089_ registers\[20\]\[48\] registers\[21\]\[48\] registers\[22\]\[48\] registers\[23\]\[48\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux4_1
XFILLER_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26705_ _11667_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ _10130_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27685_ _12214_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__clkbuf_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24897_ _10657_ VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__buf_4
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29424_ _13160_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__clkbuf_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_512 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_523 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26636_ _10814_ registers\[41\]\[40\] _11630_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__mux2_1
X_23848_ _10094_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_534 _00176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_545 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_556 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_567 _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29355_ _13068_ VGND VGND VPWR VPWR _13124_ sky130_fd_sc_hd__buf_4
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26567_ _11594_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ _10057_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_578 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_589 _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16320_ registers\[48\]\[7\] registers\[49\]\[7\] registers\[50\]\[7\] registers\[51\]\[7\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14827_ sky130_fd_sc_hd__mux4_1
X_28306_ _12541_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25518_ registers\[4\]\[25\] _10357_ _11034_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__mux2_1
XFILLER_241_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29286_ _09693_ registers\[22\]\[17\] _13080_ VGND VGND VPWR VPWR _13088_ sky130_fd_sc_hd__mux2_1
XFILLER_213_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26498_ _11557_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28237_ _12504_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__clkbuf_1
X_16251_ registers\[52\]\[5\] registers\[53\]\[5\] registers\[54\]\[5\] registers\[55\]\[5\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14760_ sky130_fd_sc_hd__mux4_1
X_25449_ _11001_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16182_ registers\[48\]\[3\] registers\[49\]\[3\] registers\[50\]\[3\] registers\[51\]\[3\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14693_ sky130_fd_sc_hd__mux4_1
X_28168_ _11792_ registers\[30\]\[30\] _12468_ VGND VGND VPWR VPWR _12469_ sky130_fd_sc_hd__mux2_1
XFILLER_166_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27119_ _11826_ registers\[38\]\[46\] _11909_ VGND VGND VPWR VPWR _11916_ sky130_fd_sc_hd__mux2_1
X_28099_ _11859_ registers\[31\]\[62\] _12363_ VGND VGND VPWR VPWR _12432_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30130_ registers\[16\]\[33\] _13004_ _13528_ VGND VGND VPWR VPWR _13532_ sky130_fd_sc_hd__mux2_1
X_19941_ _05111_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__buf_6
XFILLER_138_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30061_ registers\[16\]\[0\] _12931_ _13495_ VGND VGND VPWR VPWR _13496_ sky130_fd_sc_hd__mux2_1
X_19872_ registers\[4\]\[42\] registers\[5\]\[42\] registers\[6\]\[42\] registers\[7\]\[42\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__mux4_1
XFILLER_49_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18823_ _05501_ _05572_ _05573_ _05506_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__a22o_1
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33820_ clknet_leaf_10_CLK _01934_ VGND VGND VPWR VPWR registers\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_18754_ _05501_ _05502_ _05505_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__a22o_1
XTAP_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17705_ _14510_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__buf_4
XFILLER_82_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33751_ clknet_leaf_135_CLK _01865_ VGND VGND VPWR VPWR registers\[40\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_30963_ _13970_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_1395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18685_ registers\[32\]\[9\] registers\[33\]\[9\] registers\[34\]\[9\] registers\[35\]\[9\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__mux4_1
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32702_ clknet_leaf_290_CLK _00816_ VGND VGND VPWR VPWR registers\[57\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17636_ _15825_ _04417_ _04418_ _15828_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__a22o_1
X_33682_ clknet_leaf_128_CLK _01796_ VGND VGND VPWR VPWR registers\[41\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30894_ _13934_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35421_ clknet_leaf_480_CLK _03535_ VGND VGND VPWR VPWR registers\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_32633_ clknet_leaf_333_CLK _00747_ VGND VGND VPWR VPWR registers\[58\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17567_ _04348_ _04351_ _15963_ _15964_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__o211a_1
XFILLER_51_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19306_ _05141_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__buf_4
X_16518_ _14947_ _15018_ _15019_ _14950_ VGND VGND VPWR VPWR _15020_ sky130_fd_sc_hd__a22o_1
XFILLER_232_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35352_ clknet_leaf_44_CLK _03466_ VGND VGND VPWR VPWR registers\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_32564_ clknet_leaf_418_CLK _00678_ VGND VGND VPWR VPWR registers\[5\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17498_ registers\[4\]\[40\] registers\[5\]\[40\] registers\[6\]\[40\] registers\[7\]\[40\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _15972_ sky130_fd_sc_hd__mux4_1
XFILLER_143_1035 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34303_ clknet_leaf_273_CLK _02417_ VGND VGND VPWR VPWR registers\[32\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_31515_ _14260_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19237_ registers\[24\]\[24\] registers\[25\]\[24\] registers\[26\]\[24\] registers\[27\]\[24\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__mux4_1
X_16449_ registers\[28\]\[10\] registers\[29\]\[10\] registers\[30\]\[10\] registers\[31\]\[10\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14953_ sky130_fd_sc_hd__mux4_1
XFILLER_177_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35283_ clknet_leaf_105_CLK _03397_ VGND VGND VPWR VPWR registers\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_32495_ clknet_leaf_369_CLK _00609_ VGND VGND VPWR VPWR registers\[60\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34234_ clknet_leaf_280_CLK _02348_ VGND VGND VPWR VPWR registers\[33\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31446_ _14224_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__clkbuf_1
X_19168_ _05905_ _05908_ _05837_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__o21ba_1
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18119_ registers\[28\]\[58\] registers\[29\]\[58\] registers\[30\]\[58\] registers\[31\]\[58\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__mux4_1
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34165_ clknet_leaf_343_CLK _02279_ VGND VGND VPWR VPWR registers\[34\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31377_ registers\[7\]\[48\] net43 _14179_ VGND VGND VPWR VPWR _14188_ sky130_fd_sc_hd__mux2_1
X_19099_ _05146_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21130_ registers\[44\]\[13\] registers\[45\]\[13\] registers\[46\]\[13\] registers\[47\]\[13\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__mux4_1
X_30328_ _13635_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33116_ clknet_leaf_51_CLK _01230_ VGND VGND VPWR VPWR registers\[50\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34096_ clknet_leaf_359_CLK _02210_ VGND VGND VPWR VPWR registers\[35\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33047_ clknet_leaf_69_CLK _01161_ VGND VGND VPWR VPWR registers\[51\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_21061_ _07433_ _07747_ _07748_ _07438_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__a22o_1
XFILLER_154_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30259_ registers\[15\]\[30\] _12997_ _13599_ VGND VGND VPWR VPWR _13600_ sky130_fd_sc_hd__mux2_1
XFILLER_160_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20012_ _05141_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__buf_6
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24820_ _10639_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34998_ clknet_leaf_307_CLK _03112_ VGND VGND VPWR VPWR registers\[21\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24751_ _10603_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21963_ registers\[28\]\[36\] registers\[29\]\[36\] registers\[30\]\[36\] registers\[31\]\[36\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__mux4_1
X_33949_ clknet_leaf_22_CLK _02063_ VGND VGND VPWR VPWR registers\[37\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ _10016_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__clkbuf_8
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _07356_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__buf_6
X_27470_ _11771_ registers\[35\]\[20\] _12100_ VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__mux2_1
X_24682_ _09613_ registers\[55\]\[47\] _10558_ VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__mux2_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21894_ registers\[20\]\[34\] registers\[21\]\[34\] registers\[22\]\[34\] registers\[23\]\[34\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__mux4_1
XFILLER_82_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26421_ _11517_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__clkbuf_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35619_ clknet_leaf_466_CLK _03733_ VGND VGND VPWR VPWR registers\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_23633_ _09979_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20845_ _07440_ _07537_ _07538_ _07443_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__a22o_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29140_ _12994_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__clkbuf_1
X_26352_ _10802_ registers\[43\]\[34\] _11476_ VGND VGND VPWR VPWR _11481_ sky130_fd_sc_hd__mux2_1
X_23564_ _09942_ VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__buf_4
XFILLER_126_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20776_ _07433_ _07470_ _07471_ _07438_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__a22o_1
X_25303_ _10924_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22515_ registers\[48\]\[52\] registers\[49\]\[52\] registers\[50\]\[52\] registers\[51\]\[52\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__mux4_1
X_29071_ registers\[23\]\[6\] _12947_ _12935_ VGND VGND VPWR VPWR _12948_ sky130_fd_sc_hd__mux2_1
X_26283_ _10733_ registers\[43\]\[1\] _11443_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__mux2_1
XFILLER_167_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23495_ _09582_ registers\[19\]\[32\] _09903_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28022_ _11782_ registers\[31\]\[25\] _12386_ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__mux2_1
XFILLER_183_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25234_ _10888_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
X_22446_ _07356_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__clkbuf_8
XFILLER_167_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25165_ net52 VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__buf_4
X_22377_ registers\[0\]\[48\] registers\[1\]\[48\] registers\[2\]\[48\] registers\[3\]\[48\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__mux4_1
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24116_ _10236_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21328_ _07732_ _08007_ _08008_ _07735_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__a22o_1
X_25096_ _10801_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__clkbuf_1
X_29973_ _13449_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28924_ _12866_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21259_ _07737_ _07940_ _07941_ _07742_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__a22o_1
X_24047_ _10199_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28855_ _11805_ registers\[25\]\[36\] _12823_ VGND VGND VPWR VPWR _12830_ sky130_fd_sc_hd__mux2_1
XFILLER_77_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27806_ _12278_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__clkbuf_1
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28786_ _11736_ registers\[25\]\[3\] _12790_ VGND VGND VPWR VPWR _12794_ sky130_fd_sc_hd__mux2_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25998_ _11294_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27737_ registers\[33\]\[18\] _10342_ _12233_ VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__mux2_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24949_ _10707_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _05150_ _05229_ _05230_ _05160_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__a22o_1
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27668_ _12205_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__clkbuf_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_320 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_331 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17421_ _15892_ _15894_ _15895_ _15896_ VGND VGND VPWR VPWR _15897_ sky130_fd_sc_hd__a22o_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29407_ _09678_ registers\[21\]\[10\] _13151_ VGND VGND VPWR VPWR _13152_ sky130_fd_sc_hd__mux2_1
X_26619_ _10798_ registers\[41\]\[32\] _11619_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__mux2_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27599_ _12169_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__clkbuf_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_386 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _14510_ VGND VGND VPWR VPWR _15830_ sky130_fd_sc_hd__buf_4
XFILLER_92_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29338_ _13115_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__clkbuf_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16303_ _14588_ _14807_ _14810_ _14598_ VGND VGND VPWR VPWR _14811_ sky130_fd_sc_hd__a22o_1
XFILLER_53_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29269_ _09676_ registers\[22\]\[9\] _13069_ VGND VGND VPWR VPWR _13079_ sky130_fd_sc_hd__mux2_1
X_17283_ _15482_ _15761_ _15762_ _15485_ VGND VGND VPWR VPWR _15763_ sky130_fd_sc_hd__a22o_1
XFILLER_159_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19022_ _05127_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__buf_4
X_31300_ registers\[7\]\[11\] net3 _14146_ VGND VGND VPWR VPWR _14148_ sky130_fd_sc_hd__mux2_1
X_16234_ registers\[28\]\[4\] registers\[29\]\[4\] registers\[30\]\[4\] registers\[31\]\[4\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14744_ sky130_fd_sc_hd__mux4_1
X_32280_ clknet_leaf_8_CLK _00394_ VGND VGND VPWR VPWR registers\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31231_ _14111_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__clkbuf_1
X_16165_ _14588_ _14675_ _14676_ _14598_ VGND VGND VPWR VPWR _14677_ sky130_fd_sc_hd__a22o_1
XFILLER_126_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31162_ _14063_ VGND VGND VPWR VPWR _14075_ sky130_fd_sc_hd__buf_4
XFILLER_181_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16096_ _14515_ VGND VGND VPWR VPWR _14610_ sky130_fd_sc_hd__buf_12
XFILLER_141_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30113_ registers\[16\]\[25\] _12987_ _13517_ VGND VGND VPWR VPWR _13523_ sky130_fd_sc_hd__mux2_1
X_19924_ _06639_ _06642_ _06504_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__o21ba_1
XFILLER_130_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35970_ clknet_leaf_233_CLK _04084_ VGND VGND VPWR VPWR registers\[6\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_31093_ registers\[0\]\[41\] _13021_ _14037_ VGND VGND VPWR VPWR _14039_ sky130_fd_sc_hd__mux2_1
XFILLER_218_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30044_ _13486_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__clkbuf_1
X_34921_ clknet_leaf_454_CLK _03035_ VGND VGND VPWR VPWR registers\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_19855_ _05088_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18806_ registers\[52\]\[12\] registers\[53\]\[12\] registers\[54\]\[12\] registers\[55\]\[12\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__mux4_1
XFILLER_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34852_ clknet_leaf_472_CLK _02966_ VGND VGND VPWR VPWR registers\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19786_ registers\[60\]\[40\] registers\[61\]\[40\] registers\[62\]\[40\] registers\[63\]\[40\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__mux4_1
X_16998_ _15482_ _15483_ _15484_ _15485_ VGND VGND VPWR VPWR _15486_ sky130_fd_sc_hd__a22o_1
X_33803_ clknet_leaf_159_CLK _01917_ VGND VGND VPWR VPWR registers\[40\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18737_ _05345_ _05486_ _05489_ _05348_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__a22o_1
X_34783_ clknet_leaf_10_CLK _02897_ VGND VGND VPWR VPWR registers\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31995_ clknet_leaf_27_CLK _00167_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_1
X_33734_ clknet_leaf_248_CLK _01848_ VGND VGND VPWR VPWR registers\[41\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18668_ _05125_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__buf_6
X_30946_ _13961_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17619_ registers\[32\]\[44\] registers\[33\]\[44\] registers\[34\]\[44\] registers\[35\]\[44\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__mux4_1
XFILLER_75_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33665_ clknet_leaf_272_CLK _01779_ VGND VGND VPWR VPWR registers\[42\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30877_ _13925_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__clkbuf_1
X_18599_ registers\[24\]\[6\] registers\[25\]\[6\] registers\[26\]\[6\] registers\[27\]\[6\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__mux4_1
XFILLER_145_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35404_ clknet_leaf_150_CLK _03518_ VGND VGND VPWR VPWR registers\[15\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20630_ _07328_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__buf_4
X_32616_ clknet_leaf_436_CLK _00730_ VGND VGND VPWR VPWR registers\[58\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33596_ clknet_leaf_277_CLK _01710_ VGND VGND VPWR VPWR registers\[43\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35335_ clknet_leaf_153_CLK _03449_ VGND VGND VPWR VPWR registers\[16\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_20561_ _05040_ _07259_ _07260_ _05050_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__a22o_1
XFILLER_71_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32547_ clknet_leaf_470_CLK _00661_ VGND VGND VPWR VPWR registers\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_22300_ _07275_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__buf_4
X_35266_ clknet_leaf_223_CLK _03380_ VGND VGND VPWR VPWR registers\[17\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_20492_ registers\[56\]\[61\] registers\[57\]\[61\] registers\[58\]\[61\] registers\[59\]\[61\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__mux4_1
X_23280_ net38 VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__clkbuf_4
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32478_ clknet_leaf_50_CLK _00592_ VGND VGND VPWR VPWR registers\[60\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22231_ registers\[52\]\[44\] registers\[53\]\[44\] registers\[54\]\[44\] registers\[55\]\[44\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__mux4_1
X_34217_ clknet_leaf_431_CLK _02331_ VGND VGND VPWR VPWR registers\[33\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31429_ _14215_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35197_ clknet_leaf_191_CLK _03311_ VGND VGND VPWR VPWR registers\[18\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_246_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22162_ registers\[48\]\[42\] registers\[49\]\[42\] registers\[50\]\[42\] registers\[51\]\[42\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__mux4_1
X_34148_ clknet_leaf_56_CLK _02262_ VGND VGND VPWR VPWR registers\[34\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21113_ registers\[4\]\[12\] registers\[5\]\[12\] registers\[6\]\[12\] registers\[7\]\[12\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__mux4_1
XTAP_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26970_ _11829_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__clkbuf_1
X_22093_ _07356_ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__buf_4
XTAP_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34079_ clknet_leaf_16_CLK _02193_ VGND VGND VPWR VPWR registers\[35\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25921_ _11254_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
X_21044_ registers\[24\]\[10\] registers\[25\]\[10\] registers\[26\]\[10\] registers\[27\]\[10\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__mux4_1
XFILLER_232_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28640_ _12716_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__clkbuf_1
X_25852_ _10842_ registers\[47\]\[53\] _11214_ VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__mux2_1
X_24803_ _10630_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
X_28571_ _12680_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25783_ _10772_ registers\[47\]\[20\] _11181_ VGND VGND VPWR VPWR _11182_ sky130_fd_sc_hd__mux2_1
X_22995_ _09592_ registers\[62\]\[37\] _09578_ VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__mux2_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27522_ _11824_ registers\[35\]\[45\] _12122_ VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__mux2_1
X_24734_ _10594_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
X_21946_ _08603_ _08608_ _08405_ _08406_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__o211a_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27453_ _11755_ registers\[35\]\[12\] _12089_ VGND VGND VPWR VPWR _12092_ sky130_fd_sc_hd__mux2_1
XFILLER_203_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24665_ _09596_ registers\[55\]\[39\] _10547_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__mux2_1
XFILLER_243_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21877_ registers\[60\]\[34\] registers\[61\]\[34\] registers\[62\]\[34\] registers\[63\]\[34\]
+ _08541_ _08335_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__mux4_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26404_ _10854_ registers\[43\]\[59\] _11498_ VGND VGND VPWR VPWR _11508_ sky130_fd_sc_hd__mux2_1
XFILLER_202_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _09970_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20828_ _07519_ _07522_ _07370_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__o21ba_1
X_27384_ _12055_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__clkbuf_1
X_24596_ _09527_ registers\[55\]\[6\] _10514_ VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29123_ net16 VGND VGND VPWR VPWR _12983_ sky130_fd_sc_hd__buf_2
X_26335_ _10785_ registers\[43\]\[26\] _11465_ VGND VGND VPWR VPWR _11472_ sky130_fd_sc_hd__mux2_1
X_23547_ _09634_ registers\[19\]\[57\] _09925_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__mux2_1
XFILLER_243_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20759_ registers\[12\]\[2\] registers\[13\]\[2\] registers\[14\]\[2\] registers\[15\]\[2\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__mux4_1
X_29054_ _12936_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__clkbuf_1
X_26266_ _11435_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
X_23478_ _09565_ registers\[19\]\[24\] _09892_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__mux2_1
X_28005_ _11765_ registers\[31\]\[17\] _12375_ VGND VGND VPWR VPWR _12383_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25217_ _10879_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22429_ _07331_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__buf_4
X_26197_ _11399_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25148_ _10835_ registers\[52\]\[50\] _10836_ VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__mux2_1
XFILLER_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17970_ _04743_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_2
X_29956_ _13440_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__clkbuf_1
X_25079_ _10789_ registers\[52\]\[28\] _10773_ VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__mux2_1
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28907_ _11857_ registers\[25\]\[61\] _12789_ VGND VGND VPWR VPWR _12857_ sky130_fd_sc_hd__mux2_1
X_16921_ registers\[48\]\[24\] registers\[49\]\[24\] registers\[50\]\[24\] registers\[51\]\[24\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15411_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29887_ registers\[18\]\[46\] _13031_ _13397_ VGND VGND VPWR VPWR _13404_ sky130_fd_sc_hd__mux2_1
X_19640_ _06090_ _06365_ _06366_ _06096_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__a22o_1
XFILLER_133_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28838_ _11788_ registers\[25\]\[28\] _12812_ VGND VGND VPWR VPWR _12821_ sky130_fd_sc_hd__mux2_1
X_16852_ _14516_ VGND VGND VPWR VPWR _15344_ sky130_fd_sc_hd__buf_4
XFILLER_226_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19571_ _06296_ _06299_ _06161_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__o21ba_1
X_16783_ _14553_ VGND VGND VPWR VPWR _15277_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28769_ _12784_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_58__f_CLK clknet_5_29_0_CLK VGND VGND VPWR VPWR clknet_6_58__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_218_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18522_ registers\[8\]\[4\] registers\[9\]\[4\] registers\[10\]\[4\] registers\[11\]\[4\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__mux4_1
X_30800_ _09753_ registers\[11\]\[30\] _13884_ VGND VGND VPWR VPWR _13885_ sky130_fd_sc_hd__mux2_1
XFILLER_74_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31780_ registers\[59\]\[47\] net42 _14392_ VGND VGND VPWR VPWR _14400_ sky130_fd_sc_hd__mux2_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30731_ registers\[12\]\[62\] _13064_ _13779_ VGND VGND VPWR VPWR _13848_ sky130_fd_sc_hd__mux2_1
X_18453_ registers\[52\]\[2\] registers\[53\]\[2\] registers\[54\]\[2\] registers\[55\]\[2\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__mux4_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ registers\[44\]\[38\] registers\[45\]\[38\] registers\[46\]\[38\] registers\[47\]\[38\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15880_ sky130_fd_sc_hd__mux4_1
X_18384_ _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__buf_4
X_33450_ clknet_leaf_429_CLK _01564_ VGND VGND VPWR VPWR registers\[45\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_183 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30662_ registers\[12\]\[29\] _12995_ _13802_ VGND VGND VPWR VPWR _13812_ sky130_fd_sc_hd__mux2_1
XFILLER_221_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_194 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32401_ clknet_leaf_102_CLK _00515_ VGND VGND VPWR VPWR registers\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ registers\[36\]\[36\] registers\[37\]\[36\] registers\[38\]\[36\] registers\[39\]\[36\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15813_ sky130_fd_sc_hd__mux4_1
X_30593_ _13775_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__clkbuf_1
X_33381_ clknet_leaf_59_CLK _01495_ VGND VGND VPWR VPWR registers\[46\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35120_ clknet_leaf_377_CLK _03234_ VGND VGND VPWR VPWR registers\[1\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32332_ clknet_leaf_147_CLK _00446_ VGND VGND VPWR VPWR registers\[19\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_17266_ registers\[32\]\[34\] registers\[33\]\[34\] registers\[34\]\[34\] registers\[35\]\[34\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15746_ sky130_fd_sc_hd__mux4_1
XFILLER_201_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16217_ _14541_ VGND VGND VPWR VPWR _14727_ sky130_fd_sc_hd__buf_6
X_19005_ _05042_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__buf_4
X_32263_ clknet_leaf_236_CLK _00377_ VGND VGND VPWR VPWR registers\[39\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_35051_ clknet_leaf_401_CLK _03165_ VGND VGND VPWR VPWR registers\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17197_ _14496_ VGND VGND VPWR VPWR _15679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34002_ clknet_leaf_120_CLK _02116_ VGND VGND VPWR VPWR registers\[36\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_31214_ _14102_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__clkbuf_1
X_16148_ _14654_ _14659_ _14525_ VGND VGND VPWR VPWR _14660_ sky130_fd_sc_hd__o21ba_1
XFILLER_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32194_ clknet_leaf_460_CLK _00308_ VGND VGND VPWR VPWR registers\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31145_ _14066_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__clkbuf_1
X_16079_ _14592_ VGND VGND VPWR VPWR _14593_ sky130_fd_sc_hd__buf_6
XFILLER_103_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19907_ _06379_ _06625_ _06626_ _06382_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__a22o_1
X_35953_ clknet_leaf_378_CLK _04067_ VGND VGND VPWR VPWR registers\[6\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_31076_ registers\[0\]\[33\] _13004_ _14026_ VGND VGND VPWR VPWR _14030_ sky130_fd_sc_hd__mux2_1
XFILLER_68_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30027_ _13477_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__clkbuf_1
X_34904_ clknet_leaf_2_CLK _03018_ VGND VGND VPWR VPWR registers\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19838_ _06556_ _06559_ _06523_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35884_ clknet_leaf_391_CLK _03998_ VGND VGND VPWR VPWR registers\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34835_ clknet_leaf_103_CLK _02949_ VGND VGND VPWR VPWR registers\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xinput1 DW[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_6
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19769_ _06187_ _06491_ _06492_ _06192_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__a22o_1
XFILLER_232_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21800_ _07285_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__buf_2
XFILLER_232_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22780_ registers\[20\]\[60\] registers\[21\]\[60\] registers\[22\]\[60\] registers\[23\]\[60\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__mux4_1
X_34766_ clknet_leaf_111_CLK _02880_ VGND VGND VPWR VPWR registers\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31978_ clknet_leaf_21_CLK _00148_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_213_904 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21731_ registers\[48\]\[30\] registers\[49\]\[30\] registers\[50\]\[30\] registers\[51\]\[30\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__mux4_1
X_33717_ clknet_leaf_344_CLK _01831_ VGND VGND VPWR VPWR registers\[41\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_30929_ _13952_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__clkbuf_1
X_34697_ clknet_leaf_216_CLK _02811_ VGND VGND VPWR VPWR registers\[26\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24450_ _09519_ registers\[56\]\[2\] _10440_ VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__mux2_1
X_33648_ clknet_leaf_347_CLK _01762_ VGND VGND VPWR VPWR registers\[42\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_21662_ _08326_ _08328_ _08331_ _08332_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__a22o_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23401_ registers\[39\]\[53\] _09804_ _09851_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__mux2_1
XFILLER_196_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20613_ _07274_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__buf_12
X_24381_ _10396_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33579_ clknet_leaf_428_CLK _01693_ VGND VGND VPWR VPWR registers\[43\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21593_ _08260_ _08265_ _08062_ _08063_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__o211a_1
XFILLER_240_1449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26120_ _10840_ registers\[45\]\[52\] _11356_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23332_ _09816_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
X_35318_ clknet_leaf_310_CLK _03432_ VGND VGND VPWR VPWR registers\[16\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_20544_ _07244_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__buf_4
XFILLER_192_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26051_ _11322_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35249_ clknet_leaf_396_CLK _03363_ VGND VGND VPWR VPWR registers\[17\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_23263_ _09770_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
X_20475_ _07174_ _07177_ _05133_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__o21ba_1
X_25002_ _10737_ registers\[52\]\[3\] _10731_ VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22214_ _08766_ _08868_ _08869_ _08771_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__a22o_1
XFILLER_180_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23194_ _09727_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29810_ _13363_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__clkbuf_1
XTAP_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22145_ _08799_ _08802_ _08773_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__o21ba_1
XTAP_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29741_ _13327_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22076_ _07331_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__buf_4
X_26953_ net37 VGND VGND VPWR VPWR _11818_ sky130_fd_sc_hd__buf_4
XFILLER_59_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21027_ registers\[60\]\[10\] registers\[61\]\[10\] registers\[62\]\[10\] registers\[63\]\[10\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__mux4_1
X_25904_ _11245_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
X_29672_ registers\[1\]\[8\] _12951_ _13282_ VGND VGND VPWR VPWR _13291_ sky130_fd_sc_hd__mux2_1
X_26884_ net13 VGND VGND VPWR VPWR _11771_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28623_ _11843_ registers\[27\]\[54\] _12703_ VGND VGND VPWR VPWR _12708_ sky130_fd_sc_hd__mux2_1
X_25835_ _10825_ registers\[47\]\[45\] _11203_ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__mux2_1
XFILLER_28_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25766_ _10756_ registers\[47\]\[12\] _11170_ VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__mux2_1
X_28554_ _11774_ registers\[27\]\[21\] _12670_ VGND VGND VPWR VPWR _12672_ sky130_fd_sc_hd__mux2_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22978_ _09581_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24717_ net83 net89 VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__nand2b_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27505_ _11807_ registers\[35\]\[37\] _12111_ VGND VGND VPWR VPWR _12119_ sky130_fd_sc_hd__mux2_1
XFILLER_245_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28485_ _12635_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__clkbuf_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21929_ _08569_ _08576_ _08585_ _08592_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__or4_1
XFILLER_203_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25697_ _11135_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27436_ _11738_ registers\[35\]\[4\] _12078_ VGND VGND VPWR VPWR _12083_ sky130_fd_sc_hd__mux2_1
XFILLER_230_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _10548_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27367_ _12046_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__clkbuf_1
X_24579_ _09511_ _09654_ VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__nor2_8
XFILLER_212_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_196_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_196_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17120_ registers\[40\]\[30\] registers\[41\]\[30\] registers\[42\]\[30\] registers\[43\]\[30\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15604_ sky130_fd_sc_hd__mux4_1
X_29106_ _12971_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26318_ _10768_ registers\[43\]\[18\] _11454_ VGND VGND VPWR VPWR _11463_ sky130_fd_sc_hd__mux2_1
XFILLER_180_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27298_ _12010_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1068 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29037_ _12925_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__clkbuf_1
X_17051_ registers\[44\]\[28\] registers\[45\]\[28\] registers\[46\]\[28\] registers\[47\]\[28\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15537_ sky130_fd_sc_hd__mux4_1
X_26249_ _11426_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16002_ _14515_ VGND VGND VPWR VPWR _14516_ sky130_fd_sc_hd__buf_12
XFILLER_104_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_977 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ registers\[8\]\[53\] registers\[9\]\[53\] registers\[10\]\[53\] registers\[11\]\[53\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux4_1
X_29939_ _13431_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__clkbuf_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16904_ registers\[16\]\[23\] registers\[17\]\[23\] registers\[18\]\[23\] registers\[19\]\[23\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15395_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_120_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_120_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32950_ clknet_leaf_330_CLK _01064_ VGND VGND VPWR VPWR registers\[53\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_17884_ _04656_ _04659_ _04619_ _04620_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__o211a_1
XFILLER_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19623_ registers\[16\]\[35\] registers\[17\]\[35\] registers\[18\]\[35\] registers\[19\]\[35\]
+ _06043_ _06044_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__mux4_1
X_31901_ _09775_ registers\[49\]\[40\] _14463_ VGND VGND VPWR VPWR _14464_ sky130_fd_sc_hd__mux2_1
X_16835_ _15290_ _15326_ _15327_ _15293_ VGND VGND VPWR VPWR _15328_ sky130_fd_sc_hd__a22o_1
X_32881_ clknet_leaf_369_CLK _00995_ VGND VGND VPWR VPWR registers\[54\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_34620_ clknet_leaf_190_CLK _02734_ VGND VGND VPWR VPWR registers\[27\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_31832_ _14427_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__clkbuf_1
X_19554_ _06036_ _06282_ _06283_ _06039_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__a22o_1
X_16766_ _15260_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18505_ _05264_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34551_ clknet_leaf_312_CLK _02665_ VGND VGND VPWR VPWR registers\[28\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_19485_ _06213_ _06216_ _06180_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__o21ba_1
X_31763_ registers\[59\]\[39\] net33 _14381_ VGND VGND VPWR VPWR _14391_ sky130_fd_sc_hd__mux2_1
X_16697_ _14991_ _15191_ _15192_ _14996_ VGND VGND VPWR VPWR _15193_ sky130_fd_sc_hd__a22o_1
XFILLER_206_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33502_ clknet_leaf_32_CLK _01616_ VGND VGND VPWR VPWR registers\[44\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30714_ _13839_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__clkbuf_1
X_18436_ _05039_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__buf_4
XFILLER_22_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34482_ clknet_leaf_384_CLK _02596_ VGND VGND VPWR VPWR registers\[2\]\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31694_ registers\[59\]\[6\] net61 _14348_ VGND VGND VPWR VPWR _14355_ sky130_fd_sc_hd__mux2_1
XFILLER_146_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36221_ clknet_leaf_116_CLK _00105_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dfxtp_1
X_33433_ clknet_leaf_30_CLK _01547_ VGND VGND VPWR VPWR registers\[45\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18367_ _05064_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_187_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_187_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30645_ _13803_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36152_ clknet_leaf_336_CLK _04266_ VGND VGND VPWR VPWR registers\[49\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17318_ registers\[12\]\[35\] registers\[13\]\[35\] registers\[14\]\[35\] registers\[15\]\[35\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15797_ sky130_fd_sc_hd__mux4_1
X_33364_ clknet_leaf_124_CLK _01478_ VGND VGND VPWR VPWR registers\[46\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_30576_ _09802_ registers\[13\]\[52\] _13764_ VGND VGND VPWR VPWR _13767_ sky130_fd_sc_hd__mux2_1
X_18298_ _05051_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__buf_4
XFILLER_200_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35103_ clknet_leaf_486_CLK _03217_ VGND VGND VPWR VPWR registers\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32315_ clknet_leaf_185_CLK _00429_ VGND VGND VPWR VPWR registers\[19\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_17249_ _15482_ _15728_ _15729_ _15485_ VGND VGND VPWR VPWR _15730_ sky130_fd_sc_hd__a22o_1
X_36083_ clknet_leaf_364_CLK _04197_ VGND VGND VPWR VPWR registers\[59\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_33295_ clknet_leaf_130_CLK _01409_ VGND VGND VPWR VPWR registers\[47\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20260_ _06722_ _06968_ _06969_ _06725_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__a22o_1
XFILLER_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35034_ clknet_leaf_1_CLK _03148_ VGND VGND VPWR VPWR registers\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_32246_ clknet_leaf_336_CLK _00360_ VGND VGND VPWR VPWR registers\[39\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20191_ _06899_ _06902_ _06866_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__o21ba_1
XFILLER_157_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32177_ clknet_leaf_15_CLK _00291_ VGND VGND VPWR VPWR registers\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31128_ registers\[0\]\[58\] _13056_ _14048_ VGND VGND VPWR VPWR _14057_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_111_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_111_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23950_ _09626_ registers\[60\]\[53\] _10144_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__mux2_1
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35936_ clknet_leaf_481_CLK _04050_ VGND VGND VPWR VPWR registers\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31059_ registers\[0\]\[25\] _12987_ _14015_ VGND VGND VPWR VPWR _14021_ sky130_fd_sc_hd__mux2_1
XFILLER_57_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22901_ net62 VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35867_ clknet_leaf_476_CLK _03981_ VGND VGND VPWR VPWR registers\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_23881_ _09556_ registers\[60\]\[20\] _10111_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__mux2_1
X_25620_ registers\[48\]\[8\] _10321_ _11086_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__mux2_1
X_34818_ clknet_leaf_224_CLK _02932_ VGND VGND VPWR VPWR registers\[24\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_22832_ registers\[12\]\[62\] registers\[13\]\[62\] registers\[14\]\[62\] registers\[15\]\[62\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__mux4_1
XFILLER_72_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35798_ clknet_leaf_85_CLK _03912_ VGND VGND VPWR VPWR registers\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_908 _09685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_919 _09760_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_41__f_CLK clknet_5_20_0_CLK VGND VGND VPWR VPWR clknet_6_41__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_225_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25551_ _11057_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22763_ registers\[48\]\[60\] registers\[49\]\[60\] registers\[50\]\[60\] registers\[51\]\[60\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__mux4_1
X_34749_ clknet_leaf_182_CLK _02863_ VGND VGND VPWR VPWR registers\[25\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24502_ _09571_ registers\[56\]\[27\] _10462_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__mux2_1
X_21714_ registers\[28\]\[29\] registers\[29\]\[29\] registers\[30\]\[29\] registers\[31\]\[29\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__mux4_1
X_28270_ _12522_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__clkbuf_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25482_ registers\[4\]\[8\] _10321_ _11012_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__mux2_1
X_22694_ _09335_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27221_ _11792_ registers\[37\]\[30\] _11969_ VGND VGND VPWR VPWR _11970_ sky130_fd_sc_hd__mux2_1
X_24433_ _10431_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_178_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_178_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21645_ _08313_ _08316_ _08087_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__o21ba_1
XFILLER_21_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27152_ _11859_ registers\[38\]\[62\] _11864_ VGND VGND VPWR VPWR _11933_ sky130_fd_sc_hd__mux2_1
XFILLER_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24364_ registers\[57\]\[38\] _10384_ _10368_ VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__mux2_1
XANTENNA_50 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21576_ _08226_ _08233_ _08242_ _08249_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__or4_4
XANTENNA_61 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26103_ _10823_ registers\[45\]\[44\] _11345_ VGND VGND VPWR VPWR _11350_ sky130_fd_sc_hd__mux2_1
X_23315_ _09805_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__clkbuf_1
X_20527_ _05149_ _07226_ _07227_ _05159_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__a22o_1
XANTENNA_83 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27083_ _11790_ registers\[38\]\[29\] _11887_ VGND VGND VPWR VPWR _11897_ sky130_fd_sc_hd__mux2_1
XANTENNA_94 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24295_ net8 VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__buf_6
XFILLER_125_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26034_ _10754_ registers\[45\]\[11\] _11312_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__mux2_1
X_23246_ _09759_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
X_20458_ registers\[44\]\[60\] registers\[45\]\[60\] registers\[46\]\[60\] registers\[47\]\[60\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__mux4_1
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_350_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_350_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23177_ _09718_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XTAP_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20389_ registers\[28\]\[57\] registers\[29\]\[57\] registers\[30\]\[57\] registers\[31\]\[57\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__mux4_1
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1307 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1318 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22128_ registers\[60\]\[41\] registers\[61\]\[41\] registers\[62\]\[41\] registers\[63\]\[41\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__mux4_1
XTAP_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput190 net190 VGND VGND VPWR VPWR D2[42] sky130_fd_sc_hd__buf_2
XTAP_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27985_ _12372_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1329 _00161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29724_ _13318_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_102_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_102_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26936_ _11806_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_1
X_22059_ _08610_ _08717_ _08718_ _08613_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__a22o_1
XFILLER_82_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29655_ _13281_ VGND VGND VPWR VPWR _13282_ sky130_fd_sc_hd__buf_4
X_26867_ _11759_ registers\[3\]\[14\] _11751_ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__mux2_1
XTAP_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28606_ _11826_ registers\[27\]\[46\] _12692_ VGND VGND VPWR VPWR _12699_ sky130_fd_sc_hd__mux2_1
X_16620_ registers\[20\]\[15\] registers\[21\]\[15\] registers\[22\]\[15\] registers\[23\]\[15\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15119_ sky130_fd_sc_hd__mux4_1
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25818_ _10808_ registers\[47\]\[37\] _11192_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__mux2_1
X_26798_ _11716_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_1
X_29586_ registers\[20\]\[31\] _13000_ _13244_ VGND VGND VPWR VPWR _13246_ sky130_fd_sc_hd__mux2_1
XFILLER_16_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16551_ registers\[16\]\[13\] registers\[17\]\[13\] registers\[18\]\[13\] registers\[19\]\[13\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _15052_ sky130_fd_sc_hd__mux4_1
XFILLER_244_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25749_ _10739_ registers\[47\]\[4\] _11159_ VGND VGND VPWR VPWR _11164_ sky130_fd_sc_hd__mux2_1
X_28537_ _11757_ registers\[27\]\[13\] _12659_ VGND VGND VPWR VPWR _12663_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19270_ registers\[16\]\[25\] registers\[17\]\[25\] registers\[18\]\[25\] registers\[19\]\[25\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__mux4_1
X_16482_ _14947_ _14983_ _14984_ _14950_ VGND VGND VPWR VPWR _14985_ sky130_fd_sc_hd__a22o_1
X_28468_ _12626_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18221_ _04982_ _04985_ _14524_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__o21ba_1
XFILLER_223_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27419_ _12073_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_169_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_169_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_176_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28399_ _12590_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30430_ _09791_ registers\[14\]\[47\] _13682_ VGND VGND VPWR VPWR _13690_ sky130_fd_sc_hd__mux2_1
X_18152_ _04916_ _04919_ _04644_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__o21ba_1
XFILLER_50_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17103_ _15584_ _15587_ _15277_ _15278_ VGND VGND VPWR VPWR _15588_ sky130_fd_sc_hd__o211a_1
X_18083_ registers\[4\]\[57\] registers\[5\]\[57\] registers\[6\]\[57\] registers\[7\]\[57\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__mux4_1
XFILLER_183_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30361_ _09687_ registers\[14\]\[14\] _13649_ VGND VGND VPWR VPWR _13654_ sky130_fd_sc_hd__mux2_1
XFILLER_8_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17034_ _15482_ _15519_ _15520_ _15485_ VGND VGND VPWR VPWR _15521_ sky130_fd_sc_hd__a22o_1
X_32100_ clknet_leaf_483_CLK _00014_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33080_ clknet_leaf_337_CLK _01194_ VGND VGND VPWR VPWR registers\[51\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_30292_ registers\[15\]\[46\] _13031_ _13610_ VGND VGND VPWR VPWR _13617_ sky130_fd_sc_hd__mux2_1
XFILLER_172_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32031_ clknet_leaf_49_CLK _00209_ VGND VGND VPWR VPWR registers\[62\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_341_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_341_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _05727_ _05730_ _05494_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__o21ba_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _04705_ _04710_ _04644_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__o21ba_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33982_ clknet_leaf_269_CLK _02096_ VGND VGND VPWR VPWR registers\[37\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35721_ clknet_leaf_155_CLK _03835_ VGND VGND VPWR VPWR registers\[10\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_32933_ clknet_leaf_442_CLK _01047_ VGND VGND VPWR VPWR registers\[53\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_17867_ _14613_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__buf_2
X_19606_ registers\[56\]\[35\] registers\[57\]\[35\] registers\[58\]\[35\] registers\[59\]\[35\]
+ _06301_ _06091_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__mux4_1
X_35652_ clknet_leaf_226_CLK _03766_ VGND VGND VPWR VPWR registers\[11\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_16818_ _15307_ _15310_ _15269_ VGND VGND VPWR VPWR _15311_ sky130_fd_sc_hd__o21ba_1
XFILLER_19_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32864_ clknet_leaf_44_CLK _00978_ VGND VGND VPWR VPWR registers\[54\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_17798_ _04333_ _04572_ _04575_ _04338_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a22o_1
XFILLER_228_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34603_ clknet_leaf_452_CLK _02717_ VGND VGND VPWR VPWR registers\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_31815_ _11584_ _10512_ VGND VGND VPWR VPWR _14418_ sky130_fd_sc_hd__nand2_8
X_19537_ registers\[36\]\[33\] registers\[37\]\[33\] registers\[38\]\[33\] registers\[39\]\[33\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux4_1
XFILLER_207_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35583_ clknet_leaf_297_CLK _03697_ VGND VGND VPWR VPWR registers\[12\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_16749_ _15206_ _15242_ _15243_ _15210_ VGND VGND VPWR VPWR _15244_ sky130_fd_sc_hd__a22o_1
XFILLER_235_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32795_ clknet_leaf_54_CLK _00909_ VGND VGND VPWR VPWR registers\[55\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_34534_ clknet_leaf_455_CLK _02648_ VGND VGND VPWR VPWR registers\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31746_ _14382_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__clkbuf_1
X_19468_ registers\[44\]\[31\] registers\[45\]\[31\] registers\[46\]\[31\] registers\[47\]\[31\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__mux4_2
X_18419_ _05177_ _05180_ _05103_ _05105_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__o211a_1
XFILLER_146_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34465_ clknet_leaf_480_CLK _02579_ VGND VGND VPWR VPWR registers\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_31677_ _14345_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19399_ _06090_ _06131_ _06132_ _06096_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a22o_1
XFILLER_226_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36204_ clknet_leaf_29_CLK _00087_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dfxtp_1
X_33416_ clknet_leaf_251_CLK _01530_ VGND VGND VPWR VPWR registers\[46\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_21430_ registers\[4\]\[21\] registers\[5\]\[21\] registers\[6\]\[21\] registers\[7\]\[21\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__mux4_1
XFILLER_37_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30628_ _13794_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34396_ clknet_leaf_0_CLK _02510_ VGND VGND VPWR VPWR registers\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36135_ clknet_leaf_435_CLK _04249_ VGND VGND VPWR VPWR registers\[49\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_33347_ clknet_leaf_255_CLK _01461_ VGND VGND VPWR VPWR registers\[47\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21361_ registers\[28\]\[19\] registers\[29\]\[19\] registers\[30\]\[19\] registers\[31\]\[19\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__mux4_1
XFILLER_163_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30559_ _09784_ registers\[13\]\[44\] _13753_ VGND VGND VPWR VPWR _13758_ sky130_fd_sc_hd__mux2_1
XFILLER_159_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23100_ registers\[39\]\[4\] _09666_ _09658_ VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__mux2_1
XFILLER_174_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20312_ registers\[56\]\[55\] registers\[57\]\[55\] registers\[58\]\[55\] registers\[59\]\[55\]
+ _06987_ _06777_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__mux4_1
XFILLER_174_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput70 R1[5] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
X_24080_ _09619_ registers\[5\]\[50\] _10216_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__mux2_1
XFILLER_159_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36066_ clknet_leaf_443_CLK _04180_ VGND VGND VPWR VPWR registers\[59\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xinput81 R3[4] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
X_33278_ clknet_leaf_268_CLK _01392_ VGND VGND VPWR VPWR registers\[48\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_21292_ _07970_ _07973_ _07744_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__o21ba_1
XFILLER_200_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35017_ clknet_leaf_212_CLK _03131_ VGND VGND VPWR VPWR registers\[21\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_23031_ net44 VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__clkbuf_4
X_32229_ clknet_leaf_155_CLK _00343_ VGND VGND VPWR VPWR registers\[9\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20243_ registers\[36\]\[53\] registers\[37\]\[53\] registers\[38\]\[53\] registers\[39\]\[53\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__mux4_1
XFILLER_162_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_332_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_332_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20174_ registers\[44\]\[51\] registers\[45\]\[51\] registers\[46\]\[51\] registers\[47\]\[51\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__mux4_1
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24982_ _10724_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27770_ _12259_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23933_ _09609_ registers\[60\]\[45\] _10133_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26721_ registers\[40\]\[16\] _10338_ _11669_ VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__mux2_1
X_35919_ clknet_leaf_139_CLK _04033_ VGND VGND VPWR VPWR registers\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26652_ _10831_ registers\[41\]\[48\] _11630_ VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__mux2_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29440_ _09744_ registers\[21\]\[26\] _13162_ VGND VGND VPWR VPWR _13169_ sky130_fd_sc_hd__mux2_1
XFILLER_244_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_217_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23864_ _09540_ registers\[60\]\[12\] _10100_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__mux2_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_705 _07285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25603_ _11085_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_716 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22815_ registers\[40\]\[62\] registers\[41\]\[62\] registers\[42\]\[62\] registers\[43\]\[62\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__mux4_1
X_29371_ _13132_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__clkbuf_1
X_26583_ _10762_ registers\[41\]\[15\] _11597_ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_399_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_399_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_727 _07349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23795_ _09607_ registers\[29\]\[44\] _10061_ VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__mux2_1
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_738 _07358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_749 _07369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25534_ _11048_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_1
X_28322_ _12549_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__clkbuf_1
X_22746_ registers\[24\]\[59\] registers\[25\]\[59\] registers\[26\]\[59\] registers\[27\]\[59\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__mux4_1
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28253_ _12513_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25465_ _11011_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__buf_4
X_22677_ _09020_ _09317_ _09318_ _09024_ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__a22o_1
XFILLER_90_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_980 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27204_ _11776_ registers\[37\]\[22\] _11958_ VGND VGND VPWR VPWR _11961_ sky130_fd_sc_hd__mux2_1
X_24416_ net51 VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__buf_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21628_ registers\[60\]\[27\] registers\[61\]\[27\] registers\[62\]\[27\] registers\[63\]\[27\]
+ _08198_ _07992_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__mux4_1
X_28184_ _11809_ registers\[30\]\[38\] _12468_ VGND VGND VPWR VPWR _12477_ sky130_fd_sc_hd__mux2_1
X_25396_ _10800_ registers\[50\]\[33\] _10970_ VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__mux2_1
XFILLER_40_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27135_ _11924_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_1
X_24347_ _10373_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21559_ _08229_ _08232_ _08062_ _08063_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__o211a_1
XFILLER_165_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27066_ _11888_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24278_ registers\[57\]\[10\] _10325_ _10326_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26017_ _10737_ registers\[45\]\[3\] _11301_ VGND VGND VPWR VPWR _11305_ sky130_fd_sc_hd__mux2_1
XTAP_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23229_ registers\[9\]\[27\] _09747_ _09735_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__mux2_1
XFILLER_107_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_323_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_323_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1104 _14553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1115 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1126 _14597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1137 _14613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18770_ registers\[52\]\[11\] registers\[53\]\[11\] registers\[54\]\[11\] registers\[55\]\[11\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__mux4_1
XANTENNA_1148 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27968_ _10510_ _10014_ VGND VGND VPWR VPWR _12363_ sky130_fd_sc_hd__nand2_8
X_15982_ _14495_ VGND VGND VPWR VPWR _14496_ sky130_fd_sc_hd__buf_12
XTAP_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1159 _15713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29707_ _13309_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17721_ _04501_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_4
XFILLER_248_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26919_ net25 VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__buf_4
XTAP_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27899_ _12327_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__clkbuf_1
XTAP_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29638_ registers\[20\]\[56\] _13052_ _13266_ VGND VGND VPWR VPWR _13273_ sky130_fd_sc_hd__mux2_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ registers\[40\]\[45\] registers\[41\]\[45\] registers\[42\]\[45\] registers\[43\]\[45\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__mux4_1
XFILLER_247_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ registers\[60\]\[15\] registers\[61\]\[15\] registers\[62\]\[15\] registers\[63\]\[15\]
+ _15070_ _14864_ VGND VGND VPWR VPWR _15102_ sky130_fd_sc_hd__mux4_1
XFILLER_95_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17583_ _04362_ _04367_ _04301_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__o21ba_1
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29569_ registers\[20\]\[23\] _12983_ _13233_ VGND VGND VPWR VPWR _13237_ sky130_fd_sc_hd__mux2_1
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31600_ _14305_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__clkbuf_1
X_19322_ registers\[36\]\[27\] registers\[37\]\[27\] registers\[38\]\[27\] registers\[39\]\[27\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__mux4_1
X_16534_ registers\[56\]\[13\] registers\[57\]\[13\] registers\[58\]\[13\] registers\[59\]\[13\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _15035_ sky130_fd_sc_hd__mux4_1
XFILLER_1_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32580_ clknet_leaf_231_CLK _00694_ VGND VGND VPWR VPWR registers\[5\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31531_ _09813_ registers\[6\]\[57\] _14261_ VGND VGND VPWR VPWR _14269_ sky130_fd_sc_hd__mux2_1
X_19253_ registers\[56\]\[25\] registers\[57\]\[25\] registers\[58\]\[25\] registers\[59\]\[25\]
+ _05958_ _05748_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__mux4_1
X_16465_ _14964_ _14967_ _14926_ VGND VGND VPWR VPWR _14968_ sky130_fd_sc_hd__o21ba_1
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18204_ _14511_ _04968_ _04969_ _14517_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__a22o_1
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34250_ clknet_leaf_156_CLK _02364_ VGND VGND VPWR VPWR registers\[33\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16396_ _14863_ _14899_ _14900_ _14867_ VGND VGND VPWR VPWR _14901_ sky130_fd_sc_hd__a22o_1
X_31462_ _09740_ registers\[6\]\[24\] _14228_ VGND VGND VPWR VPWR _14233_ sky130_fd_sc_hd__mux2_1
X_19184_ registers\[36\]\[23\] registers\[37\]\[23\] registers\[38\]\[23\] registers\[39\]\[23\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__mux4_1
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33201_ clknet_leaf_378_CLK _01315_ VGND VGND VPWR VPWR registers\[4\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_18135_ registers\[60\]\[59\] registers\[61\]\[59\] registers\[62\]\[59\] registers\[63\]\[59\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__mux4_1
X_30413_ _09773_ registers\[14\]\[39\] _13671_ VGND VGND VPWR VPWR _13681_ sky130_fd_sc_hd__mux2_1
X_34181_ clknet_leaf_246_CLK _02295_ VGND VGND VPWR VPWR registers\[34\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_31393_ _14196_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33132_ clknet_leaf_379_CLK _01246_ VGND VGND VPWR VPWR registers\[50\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_18066_ registers\[32\]\[57\] registers\[33\]\[57\] registers\[34\]\[57\] registers\[35\]\[57\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__mux4_1
X_30344_ _09670_ registers\[14\]\[6\] _13638_ VGND VGND VPWR VPWR _13645_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17017_ registers\[32\]\[27\] registers\[33\]\[27\] registers\[34\]\[27\] registers\[35\]\[27\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15504_ sky130_fd_sc_hd__mux4_1
Xclkbuf_6_5__f_CLK clknet_5_2_0_CLK VGND VGND VPWR VPWR clknet_6_5__leaf_CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_314_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_314_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30275_ registers\[15\]\[38\] _13014_ _13599_ VGND VGND VPWR VPWR _13608_ sky130_fd_sc_hd__mux2_1
X_33063_ clknet_leaf_434_CLK _01177_ VGND VGND VPWR VPWR registers\[51\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32014_ clknet_leaf_178_CLK _00192_ VGND VGND VPWR VPWR registers\[62\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18968_ _05122_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__buf_4
XANTENNA_1660 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1671 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_224_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17919_ _04548_ _04692_ _04693_ _04552_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__a22o_1
XANTENNA_1682 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33965_ clknet_leaf_325_CLK _02079_ VGND VGND VPWR VPWR registers\[37\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1693 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18899_ _05643_ _05646_ _05475_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__o21ba_1
X_35704_ clknet_leaf_317_CLK _03818_ VGND VGND VPWR VPWR registers\[10\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_20930_ registers\[4\]\[7\] registers\[5\]\[7\] registers\[6\]\[7\] registers\[7\]\[7\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__mux4_1
X_32916_ clknet_leaf_63_CLK _01030_ VGND VGND VPWR VPWR registers\[53\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33896_ clknet_leaf_434_CLK _02010_ VGND VGND VPWR VPWR registers\[38\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35635_ clknet_leaf_354_CLK _03749_ VGND VGND VPWR VPWR registers\[11\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20861_ _07355_ _07553_ _07554_ _07367_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__a22o_1
X_32847_ clknet_leaf_173_CLK _00961_ VGND VGND VPWR VPWR registers\[54\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22600_ registers\[20\]\[54\] registers\[21\]\[54\] registers\[22\]\[54\] registers\[23\]\[54\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__mux4_1
XFILLER_179_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23580_ _09951_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
X_35566_ clknet_leaf_392_CLK _03680_ VGND VGND VPWR VPWR registers\[12\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_32778_ clknet_leaf_177_CLK _00892_ VGND VGND VPWR VPWR registers\[56\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_20792_ _07358_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__buf_4
XFILLER_241_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22531_ _07361_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__buf_6
X_34517_ clknet_leaf_96_CLK _02631_ VGND VGND VPWR VPWR registers\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31729_ _14373_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__clkbuf_1
X_35497_ clknet_leaf_398_CLK _03611_ VGND VGND VPWR VPWR registers\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25250_ _10896_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__clkbuf_1
X_34448_ clknet_leaf_110_CLK _02562_ VGND VGND VPWR VPWR registers\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_22462_ _07315_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__buf_4
XFILLER_183_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24201_ _09605_ registers\[58\]\[43\] _10277_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__mux2_1
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21413_ registers\[32\]\[21\] registers\[33\]\[21\] registers\[34\]\[21\] registers\[35\]\[21\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__mux4_1
X_25181_ _10858_ registers\[52\]\[61\] _10730_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__mux2_1
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34379_ clknet_leaf_143_CLK _02493_ VGND VGND VPWR VPWR registers\[31\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_22393_ _09043_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
X_36118_ clknet_leaf_68_CLK _04232_ VGND VGND VPWR VPWR registers\[49\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_24132_ _09535_ registers\[58\]\[10\] _10244_ VGND VGND VPWR VPWR _10245_ sky130_fd_sc_hd__mux2_1
X_21344_ registers\[56\]\[19\] registers\[57\]\[19\] registers\[58\]\[19\] registers\[59\]\[19\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__mux4_1
XFILLER_102_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36049_ clknet_leaf_73_CLK _04163_ VGND VGND VPWR VPWR registers\[59\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_24063_ _09603_ registers\[5\]\[42\] _10205_ VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__mux2_1
X_28940_ registers\[24\]\[12\] _10330_ _12872_ VGND VGND VPWR VPWR _12875_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_305_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_305_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21275_ registers\[60\]\[17\] registers\[61\]\[17\] registers\[62\]\[17\] registers\[63\]\[17\]
+ _07855_ _07649_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__mux4_1
XFILLER_11_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23014_ _09605_ registers\[62\]\[43\] _09599_ VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__mux2_1
XFILLER_85_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20226_ _06722_ _06935_ _06936_ _06725_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__a22o_1
X_28871_ _12838_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27822_ _12286_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20157_ registers\[16\]\[50\] registers\[17\]\[50\] registers\[18\]\[50\] registers\[19\]\[50\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__mux4_1
XFILLER_213_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24965_ _09624_ registers\[53\]\[52\] _10713_ VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__mux2_1
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27753_ _12250_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20088_ registers\[28\]\[48\] registers\[29\]\[48\] registers\[30\]\[48\] registers\[31\]\[48\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux4_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26704_ registers\[40\]\[8\] _10321_ _11658_ VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__mux2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _09592_ registers\[60\]\[37\] _10122_ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__mux2_1
X_27684_ registers\[34\]\[57\] _10424_ _12206_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__mux2_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24896_ _10679_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29423_ _09695_ registers\[21\]\[18\] _13151_ VGND VGND VPWR VPWR _13160_ sky130_fd_sc_hd__mux2_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26635_ _11585_ VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__buf_4
X_23847_ _09523_ registers\[60\]\[4\] _10089_ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__mux2_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_513 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_524 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_535 _00176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_546 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_557 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29354_ _13123_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__clkbuf_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26566_ _10745_ registers\[41\]\[7\] _11586_ VGND VGND VPWR VPWR _11594_ sky130_fd_sc_hd__mux2_1
XFILLER_232_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_568 _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23778_ _09590_ registers\[29\]\[36\] _10050_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__mux2_1
XFILLER_220_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_579 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_241_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28305_ registers\[2\]\[31\] _10370_ _12539_ VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__mux2_1
XFILLER_41_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22729_ registers\[36\]\[59\] registers\[37\]\[59\] registers\[38\]\[59\] registers\[39\]\[59\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__mux4_1
X_25517_ _11039_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__clkbuf_1
X_29285_ _13087_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26497_ _10812_ registers\[42\]\[39\] _11547_ VGND VGND VPWR VPWR _11557_ sky130_fd_sc_hd__mux2_1
XFILLER_198_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16250_ registers\[60\]\[5\] registers\[61\]\[5\] registers\[62\]\[5\] registers\[63\]\[5\]
+ _14727_ _14544_ VGND VGND VPWR VPWR _14759_ sky130_fd_sc_hd__mux4_1
X_28236_ _11861_ registers\[30\]\[63\] _12434_ VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__mux2_1
X_25448_ _10852_ registers\[50\]\[58\] _10992_ VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__mux2_1
XFILLER_167_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16181_ registers\[56\]\[3\] registers\[57\]\[3\] registers\[58\]\[3\] registers\[59\]\[3\]
+ _14530_ _14532_ VGND VGND VPWR VPWR _14692_ sky130_fd_sc_hd__mux4_1
X_28167_ _12434_ VGND VGND VPWR VPWR _12468_ sky130_fd_sc_hd__buf_4
X_25379_ _10783_ registers\[50\]\[25\] _10959_ VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27118_ _11915_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__clkbuf_1
X_28098_ _12431_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19940_ _06655_ _06658_ _06523_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__o21ba_1
X_27049_ _11879_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__clkbuf_1
X_30060_ _13494_ VGND VGND VPWR VPWR _13495_ sky130_fd_sc_hd__buf_6
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19871_ registers\[12\]\[42\] registers\[13\]\[42\] registers\[14\]\[42\] registers\[15\]\[42\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__mux4_1
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18822_ registers\[20\]\[12\] registers\[21\]\[12\] registers\[22\]\[12\] registers\[23\]\[12\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__mux4_1
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18753_ _05159_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__buf_4
XTAP_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17704_ _04481_ _04482_ _04483_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__a22o_1
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33750_ clknet_leaf_128_CLK _01864_ VGND VGND VPWR VPWR registers\[40\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30962_ registers\[10\]\[43\] _13025_ _13966_ VGND VGND VPWR VPWR _13970_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18684_ _05069_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__buf_4
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32701_ clknet_leaf_290_CLK _00815_ VGND VGND VPWR VPWR registers\[57\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17635_ registers\[0\]\[44\] registers\[1\]\[44\] registers\[2\]\[44\] registers\[3\]\[44\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__mux4_1
X_33681_ clknet_leaf_130_CLK _01795_ VGND VGND VPWR VPWR registers\[41\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30893_ registers\[10\]\[10\] _12955_ _13933_ VGND VGND VPWR VPWR _13934_ sky130_fd_sc_hd__mux2_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35420_ clknet_leaf_477_CLK _03534_ VGND VGND VPWR VPWR registers\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_32632_ clknet_leaf_333_CLK _00746_ VGND VGND VPWR VPWR registers\[58\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17566_ _15892_ _04349_ _04350_ _15896_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__a22o_1
XFILLER_223_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19305_ registers\[24\]\[26\] registers\[25\]\[26\] registers\[26\]\[26\] registers\[27\]\[26\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__mux4_1
X_35351_ clknet_leaf_83_CLK _03465_ VGND VGND VPWR VPWR registers\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16517_ registers\[16\]\[12\] registers\[17\]\[12\] registers\[18\]\[12\] registers\[19\]\[12\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _15019_ sky130_fd_sc_hd__mux4_1
XFILLER_182_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32563_ clknet_leaf_380_CLK _00677_ VGND VGND VPWR VPWR registers\[5\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17497_ registers\[12\]\[40\] registers\[13\]\[40\] registers\[14\]\[40\] registers\[15\]\[40\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15971_ sky130_fd_sc_hd__mux4_1
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34302_ clknet_leaf_275_CLK _02416_ VGND VGND VPWR VPWR registers\[32\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31514_ _09795_ registers\[6\]\[49\] _14250_ VGND VGND VPWR VPWR _14260_ sky130_fd_sc_hd__mux2_1
X_19236_ _05113_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__buf_4
X_35282_ clknet_leaf_101_CLK _03396_ VGND VGND VPWR VPWR registers\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16448_ _14600_ VGND VGND VPWR VPWR _14952_ sky130_fd_sc_hd__clkbuf_4
X_32494_ clknet_leaf_370_CLK _00608_ VGND VGND VPWR VPWR registers\[60\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34233_ clknet_leaf_340_CLK _02347_ VGND VGND VPWR VPWR registers\[33\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31445_ _09691_ registers\[6\]\[16\] _14217_ VGND VGND VPWR VPWR _14224_ sky130_fd_sc_hd__mux2_1
X_19167_ _05693_ _05906_ _05907_ _05696_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a22o_1
X_16379_ _14881_ _14884_ _14614_ VGND VGND VPWR VPWR _14885_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_91_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18118_ _04632_ _04885_ _04886_ _04635_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__a22o_1
XFILLER_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34164_ clknet_leaf_349_CLK _02278_ VGND VGND VPWR VPWR registers\[34\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_31376_ _14187_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__clkbuf_1
X_19098_ registers\[16\]\[20\] registers\[17\]\[20\] registers\[18\]\[20\] registers\[19\]\[20\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__mux4_1
XFILLER_219_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33115_ clknet_leaf_35_CLK _01229_ VGND VGND VPWR VPWR registers\[50\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_18049_ registers\[8\]\[56\] registers\[9\]\[56\] registers\[10\]\[56\] registers\[11\]\[56\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__mux4_1
X_30327_ registers\[15\]\[63\] _13066_ _13565_ VGND VGND VPWR VPWR _13635_ sky130_fd_sc_hd__mux2_1
XFILLER_219_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34095_ clknet_leaf_355_CLK _02209_ VGND VGND VPWR VPWR registers\[35\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33046_ clknet_leaf_68_CLK _01160_ VGND VGND VPWR VPWR registers\[51\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_21060_ registers\[32\]\[11\] registers\[33\]\[11\] registers\[34\]\[11\] registers\[35\]\[11\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__mux4_1
X_30258_ _13565_ VGND VGND VPWR VPWR _13599_ sky130_fd_sc_hd__buf_6
XFILLER_87_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20011_ registers\[24\]\[46\] registers\[25\]\[46\] registers\[26\]\[46\] registers\[27\]\[46\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__mux4_1
XFILLER_101_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30189_ _13562_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34997_ clknet_leaf_384_CLK _03111_ VGND VGND VPWR VPWR registers\[21\]\[39\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1490 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24750_ _09544_ registers\[54\]\[14\] _10598_ VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__mux2_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21962_ _08418_ _08621_ _08624_ _08421_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__a22o_1
X_33948_ clknet_leaf_23_CLK _02062_ VGND VGND VPWR VPWR registers\[37\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23701_ _10014_ _10015_ VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__nand2_8
XFILLER_215_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20913_ registers\[44\]\[7\] registers\[45\]\[7\] registers\[46\]\[7\] registers\[47\]\[7\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__mux4_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24681_ _10565_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
X_33879_ clknet_leaf_117_CLK _01993_ VGND VGND VPWR VPWR registers\[38\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_21893_ registers\[28\]\[34\] registers\[29\]\[34\] registers\[30\]\[34\] registers\[31\]\[34\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__mux4_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26420_ _10735_ registers\[42\]\[2\] _11514_ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__mux2_1
X_23632_ registers\[61\]\[32\] _09758_ _09976_ VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__mux2_1
X_35618_ clknet_leaf_466_CLK _03732_ VGND VGND VPWR VPWR registers\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20844_ registers\[36\]\[5\] registers\[37\]\[5\] registers\[38\]\[5\] registers\[39\]\[5\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__mux4_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_20_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_20_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_202_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26351_ _11480_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__clkbuf_1
X_23563_ _09940_ _09941_ VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__nor2_8
X_35549_ clknet_leaf_480_CLK _03663_ VGND VGND VPWR VPWR registers\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_20775_ registers\[32\]\[3\] registers\[33\]\[3\] registers\[34\]\[3\] registers\[35\]\[3\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__mux4_1
XFILLER_39_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25302_ _10842_ registers\[51\]\[53\] _10920_ VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__mux2_1
XFILLER_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22514_ registers\[56\]\[52\] registers\[57\]\[52\] registers\[58\]\[52\] registers\[59\]\[52\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__mux4_1
X_26282_ _11444_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
X_29070_ net61 VGND VGND VPWR VPWR _12947_ sky130_fd_sc_hd__clkbuf_4
XFILLER_11_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23494_ _09905_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28021_ _12391_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__clkbuf_1
X_25233_ _10772_ registers\[51\]\[20\] _10887_ VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__mux2_1
X_22445_ registers\[8\]\[50\] registers\[9\]\[50\] registers\[10\]\[50\] registers\[11\]\[50\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__mux4_1
XFILLER_210_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_82_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25164_ _10847_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__clkbuf_1
X_22376_ registers\[8\]\[48\] registers\[9\]\[48\] registers\[10\]\[48\] registers\[11\]\[48\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__mux4_1
XFILLER_100_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24115_ _09519_ registers\[58\]\[2\] _10233_ VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__mux2_1
XFILLER_135_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21327_ registers\[16\]\[18\] registers\[17\]\[18\] registers\[18\]\[18\] registers\[19\]\[18\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__mux4_1
XFILLER_191_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25095_ _10800_ registers\[52\]\[33\] _10794_ VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__mux2_1
X_29972_ registers\[17\]\[22\] _12981_ _13446_ VGND VGND VPWR VPWR _13449_ sky130_fd_sc_hd__mux2_1
X_28923_ registers\[24\]\[4\] _10313_ _12861_ VGND VGND VPWR VPWR _12866_ sky130_fd_sc_hd__mux2_1
X_24046_ _09586_ registers\[5\]\[34\] _10194_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__mux2_1
XFILLER_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21258_ registers\[20\]\[16\] registers\[21\]\[16\] registers\[22\]\[16\] registers\[23\]\[16\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__mux4_1
XFILLER_104_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20209_ registers\[44\]\[52\] registers\[45\]\[52\] registers\[46\]\[52\] registers\[47\]\[52\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__mux4_1
XFILLER_150_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28854_ _12829_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21189_ _07737_ _07872_ _07873_ _07742_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__a22o_1
XFILLER_78_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27805_ registers\[33\]\[50\] _10409_ _12277_ VGND VGND VPWR VPWR _12278_ sky130_fd_sc_hd__mux2_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28785_ _12793_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__clkbuf_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25997_ _10852_ registers\[46\]\[58\] _11285_ VGND VGND VPWR VPWR _11294_ sky130_fd_sc_hd__mux2_1
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27736_ _12241_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__clkbuf_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24948_ _09607_ registers\[53\]\[44\] _10702_ VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__mux2_1
XFILLER_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27667_ registers\[34\]\[49\] _10407_ _12195_ VGND VGND VPWR VPWR _12205_ sky130_fd_sc_hd__mux2_1
XANTENNA_310 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24879_ _09538_ registers\[53\]\[11\] _10669_ VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__mux2_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_332 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29406_ _13139_ VGND VGND VPWR VPWR _13151_ sky130_fd_sc_hd__buf_4
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17420_ _14516_ VGND VGND VPWR VPWR _15896_ sky130_fd_sc_hd__clkbuf_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_343 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26618_ _11621_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_354 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27598_ registers\[34\]\[16\] _10338_ _12162_ VGND VGND VPWR VPWR _12169_ sky130_fd_sc_hd__mux2_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_376 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29337_ _09778_ registers\[22\]\[41\] _13113_ VGND VGND VPWR VPWR _13115_ sky130_fd_sc_hd__mux2_1
X_17351_ _15825_ _15826_ _15827_ _15828_ VGND VGND VPWR VPWR _15829_ sky130_fd_sc_hd__a22o_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26549_ net85 net84 _09654_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__nor3_4
XANTENNA_398 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16302_ registers\[16\]\[6\] registers\[17\]\[6\] registers\[18\]\[6\] registers\[19\]\[6\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14810_ sky130_fd_sc_hd__mux4_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29268_ _13078_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17282_ registers\[0\]\[34\] registers\[1\]\[34\] registers\[2\]\[34\] registers\[3\]\[34\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15762_ sky130_fd_sc_hd__mux4_1
XFILLER_158_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19021_ _05125_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__buf_6
X_28219_ _12495_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__clkbuf_1
X_16233_ _14588_ _14741_ _14742_ _14598_ VGND VGND VPWR VPWR _14743_ sky130_fd_sc_hd__a22o_1
XFILLER_174_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29199_ _13034_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_73_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_73_CLK sky130_fd_sc_hd__clkbuf_16
X_31230_ registers\[8\]\[42\] net37 _14108_ VGND VGND VPWR VPWR _14111_ sky130_fd_sc_hd__mux2_1
X_16164_ registers\[16\]\[2\] registers\[17\]\[2\] registers\[18\]\[2\] registers\[19\]\[2\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14676_ sky130_fd_sc_hd__mux4_1
XFILLER_166_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_18__f_CLK clknet_5_9_0_CLK VGND VGND VPWR VPWR clknet_6_18__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_220_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16095_ registers\[20\]\[0\] registers\[21\]\[0\] registers\[22\]\[0\] registers\[23\]\[0\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14609_ sky130_fd_sc_hd__mux4_1
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31161_ _14074_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19923_ _06576_ _06640_ _06641_ _06579_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__a22o_1
XFILLER_29_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30112_ _13522_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_218_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31092_ _14038_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30043_ registers\[17\]\[56\] _13052_ _13479_ VGND VGND VPWR VPWR _13486_ sky130_fd_sc_hd__mux2_1
X_34920_ clknet_leaf_457_CLK _03034_ VGND VGND VPWR VPWR registers\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_19854_ _06569_ _06572_ _06573_ _06574_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__a22o_1
XFILLER_116_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18805_ registers\[60\]\[12\] registers\[61\]\[12\] registers\[62\]\[12\] registers\[63\]\[12\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__mux4_1
X_34851_ clknet_leaf_473_CLK _02965_ VGND VGND VPWR VPWR registers\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19785_ _06433_ _06506_ _06507_ _06439_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__a22o_1
XFILLER_110_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16997_ _14567_ VGND VGND VPWR VPWR _15485_ sky130_fd_sc_hd__buf_4
XFILLER_37_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33802_ clknet_leaf_161_CLK _01916_ VGND VGND VPWR VPWR registers\[40\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18736_ registers\[0\]\[10\] registers\[1\]\[10\] registers\[2\]\[10\] registers\[3\]\[10\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__mux4_1
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34782_ clknet_leaf_3_CLK _02896_ VGND VGND VPWR VPWR registers\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31994_ clknet_leaf_23_CLK _00166_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_1
XFILLER_236_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33733_ clknet_leaf_250_CLK _01847_ VGND VGND VPWR VPWR registers\[41\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18667_ registers\[12\]\[8\] registers\[13\]\[8\] registers\[14\]\[8\] registers\[15\]\[8\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__mux4_1
X_30945_ registers\[10\]\[35\] _13008_ _13955_ VGND VGND VPWR VPWR _13961_ sky130_fd_sc_hd__mux2_1
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17618_ registers\[40\]\[44\] registers\[41\]\[44\] registers\[42\]\[44\] registers\[43\]\[44\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__mux4_1
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33664_ clknet_leaf_272_CLK _01778_ VGND VGND VPWR VPWR registers\[42\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30876_ registers\[10\]\[2\] _12939_ _13922_ VGND VGND VPWR VPWR _13925_ sky130_fd_sc_hd__mux2_1
X_18598_ _05349_ _05354_ _05134_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__o21ba_1
XFILLER_149_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35403_ clknet_leaf_150_CLK _03517_ VGND VGND VPWR VPWR registers\[15\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_32615_ clknet_leaf_437_CLK _00729_ VGND VGND VPWR VPWR registers\[58\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17549_ _14493_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__buf_4
X_33595_ clknet_leaf_278_CLK _01709_ VGND VGND VPWR VPWR registers\[43\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_35334_ clknet_leaf_154_CLK _03448_ VGND VGND VPWR VPWR registers\[16\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20560_ registers\[0\]\[63\] registers\[1\]\[63\] registers\[2\]\[63\] registers\[3\]\[63\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__mux4_1
XFILLER_225_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32546_ clknet_leaf_470_CLK _00660_ VGND VGND VPWR VPWR registers\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19219_ _05078_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__buf_6
X_35265_ clknet_leaf_221_CLK _03379_ VGND VGND VPWR VPWR registers\[17\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_20491_ _07189_ _07192_ _05073_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32477_ clknet_leaf_57_CLK _00591_ VGND VGND VPWR VPWR registers\[60\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_64_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_64_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22230_ registers\[60\]\[44\] registers\[61\]\[44\] registers\[62\]\[44\] registers\[63\]\[44\]
+ _08884_ _08678_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__mux4_1
XFILLER_118_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34216_ clknet_leaf_430_CLK _02330_ VGND VGND VPWR VPWR registers\[33\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31428_ _09674_ registers\[6\]\[8\] _14206_ VGND VGND VPWR VPWR _14215_ sky130_fd_sc_hd__mux2_1
X_35196_ clknet_leaf_190_CLK _03310_ VGND VGND VPWR VPWR registers\[18\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22161_ registers\[56\]\[42\] registers\[57\]\[42\] registers\[58\]\[42\] registers\[59\]\[42\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__mux4_1
X_34147_ clknet_leaf_49_CLK _02261_ VGND VGND VPWR VPWR registers\[34\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31359_ _14178_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21112_ registers\[12\]\[12\] registers\[13\]\[12\] registers\[14\]\[12\] registers\[15\]\[12\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__mux4_1
XTAP_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34078_ clknet_leaf_22_CLK _02192_ VGND VGND VPWR VPWR registers\[35\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_22092_ registers\[8\]\[40\] registers\[9\]\[40\] registers\[10\]\[40\] registers\[11\]\[40\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__mux4_1
XTAP_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33029_ clknet_leaf_270_CLK _01143_ VGND VGND VPWR VPWR registers\[52\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_25920_ _10775_ registers\[46\]\[21\] _11252_ VGND VGND VPWR VPWR _11254_ sky130_fd_sc_hd__mux2_1
X_21043_ _07372_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_236_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25851_ _11217_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24802_ _09596_ registers\[54\]\[39\] _10620_ VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__mux2_1
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28570_ _11790_ registers\[27\]\[29\] _12670_ VGND VGND VPWR VPWR _12680_ sky130_fd_sc_hd__mux2_1
XFILLER_132_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25782_ _11158_ VGND VGND VPWR VPWR _11181_ sky130_fd_sc_hd__buf_4
X_22994_ net31 VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__buf_4
XFILLER_228_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27521_ _12127_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24733_ _09527_ registers\[54\]\[6\] _10587_ VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__mux2_1
XFILLER_131_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21945_ _08334_ _08604_ _08607_ _08338_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__a22o_1
XFILLER_83_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27452_ _12091_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__clkbuf_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _10556_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _07326_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__buf_6
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26403_ _11507_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__clkbuf_1
X_23615_ registers\[61\]\[24\] _09740_ _09965_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__mux2_1
XFILLER_70_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20827_ _07355_ _07520_ _07521_ _07367_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__a22o_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24595_ _10520_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
X_27383_ registers\[36\]\[43\] _10395_ _12051_ VGND VGND VPWR VPWR _12055_ sky130_fd_sc_hd__mux2_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29122_ _12982_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23546_ _09932_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26334_ _11471_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20758_ _07343_ _07453_ _07454_ _07353_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__a22o_1
XFILLER_195_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26265_ _10850_ registers\[44\]\[57\] _11427_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__mux2_1
X_29053_ registers\[23\]\[0\] _12931_ _12935_ VGND VGND VPWR VPWR _12936_ sky130_fd_sc_hd__mux2_1
X_23477_ _09896_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20689_ _07316_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_55_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_55_CLK sky130_fd_sc_hd__clkbuf_16
X_25216_ _10756_ registers\[51\]\[12\] _10876_ VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__mux2_1
X_28004_ _12382_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22428_ _08805_ _09075_ _09076_ _08810_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__a22o_1
X_26196_ _10781_ registers\[44\]\[24\] _11394_ VGND VGND VPWR VPWR _11399_ sky130_fd_sc_hd__mux2_1
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25147_ _10730_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__buf_6
X_22359_ _08812_ _09008_ _09009_ _08815_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__a22o_1
XFILLER_136_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29955_ registers\[17\]\[14\] _12964_ _13435_ VGND VGND VPWR VPWR _13440_ sky130_fd_sc_hd__mux2_1
X_25078_ net21 VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__buf_2
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28906_ _12856_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__clkbuf_1
X_24029_ _09569_ registers\[5\]\[26\] _10183_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__mux2_1
X_16920_ registers\[56\]\[24\] registers\[57\]\[24\] registers\[58\]\[24\] registers\[59\]\[24\]
+ _15409_ _15199_ VGND VGND VPWR VPWR _15410_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29886_ _13403_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28837_ _12820_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__clkbuf_1
X_16851_ registers\[36\]\[22\] registers\[37\]\[22\] registers\[38\]\[22\] registers\[39\]\[22\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15343_ sky130_fd_sc_hd__mux4_1
XFILLER_24_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19570_ _06233_ _06297_ _06298_ _06236_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__a22o_1
XFILLER_77_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28768_ _11853_ registers\[26\]\[59\] _12774_ VGND VGND VPWR VPWR _12784_ sky130_fd_sc_hd__mux2_1
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16782_ _15206_ _15274_ _15275_ _15210_ VGND VGND VPWR VPWR _15276_ sky130_fd_sc_hd__a22o_1
XFILLER_93_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18521_ _05275_ _05279_ _05103_ _05105_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__o211a_1
X_27719_ _12232_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__clkbuf_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28699_ _11784_ registers\[26\]\[26\] _12741_ VGND VGND VPWR VPWR _12748_ sky130_fd_sc_hd__mux2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30730_ _13847_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__clkbuf_1
X_18452_ registers\[60\]\[2\] registers\[61\]\[2\] registers\[62\]\[2\] registers\[63\]\[2\]
+ _05091_ _05093_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux4_1
XFILLER_146_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17403_ _15677_ _15877_ _15878_ _15682_ VGND VGND VPWR VPWR _15879_ sky130_fd_sc_hd__a22o_1
XANTENNA_173 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _05048_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__buf_12
X_30661_ _13811_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_184 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32400_ clknet_leaf_114_CLK _00514_ VGND VGND VPWR VPWR registers\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ registers\[44\]\[36\] registers\[45\]\[36\] registers\[46\]\[36\] registers\[47\]\[36\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15812_ sky130_fd_sc_hd__mux4_1
X_33380_ clknet_leaf_62_CLK _01494_ VGND VGND VPWR VPWR registers\[46\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_30592_ _09819_ registers\[13\]\[60\] _13708_ VGND VGND VPWR VPWR _13775_ sky130_fd_sc_hd__mux2_1
XFILLER_222_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32331_ clknet_leaf_149_CLK _00445_ VGND VGND VPWR VPWR registers\[19\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17265_ registers\[40\]\[34\] registers\[41\]\[34\] registers\[42\]\[34\] registers\[43\]\[34\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15745_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_46_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_46_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19004_ registers\[56\]\[18\] registers\[57\]\[18\] registers\[58\]\[18\] registers\[59\]\[18\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__mux4_1
X_16216_ _14528_ _14724_ _14725_ _14537_ VGND VGND VPWR VPWR _14726_ sky130_fd_sc_hd__a22o_1
X_35050_ clknet_leaf_405_CLK _03164_ VGND VGND VPWR VPWR registers\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_32262_ clknet_leaf_253_CLK _00376_ VGND VGND VPWR VPWR registers\[39\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17196_ _14493_ VGND VGND VPWR VPWR _15678_ sky130_fd_sc_hd__buf_4
X_34001_ clknet_leaf_134_CLK _02115_ VGND VGND VPWR VPWR registers\[36\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31213_ registers\[8\]\[34\] net28 _14097_ VGND VGND VPWR VPWR _14102_ sky130_fd_sc_hd__mux2_1
X_16147_ _14655_ _14656_ _14657_ _14658_ VGND VGND VPWR VPWR _14659_ sky130_fd_sc_hd__a22o_1
XFILLER_182_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32193_ clknet_leaf_434_CLK _00307_ VGND VGND VPWR VPWR registers\[39\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31144_ registers\[8\]\[1\] net12 _14064_ VGND VGND VPWR VPWR _14066_ sky130_fd_sc_hd__mux2_1
XFILLER_143_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16078_ _14529_ VGND VGND VPWR VPWR _14592_ sky130_fd_sc_hd__buf_12
XFILLER_115_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19906_ registers\[4\]\[43\] registers\[5\]\[43\] registers\[6\]\[43\] registers\[7\]\[43\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__mux4_1
X_31075_ _14029_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__clkbuf_1
X_35952_ clknet_leaf_374_CLK _04066_ VGND VGND VPWR VPWR registers\[6\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34903_ clknet_leaf_99_CLK _03017_ VGND VGND VPWR VPWR registers\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_30026_ registers\[17\]\[48\] _13035_ _13468_ VGND VGND VPWR VPWR _13477_ sky130_fd_sc_hd__mux2_1
X_19837_ _06379_ _06557_ _06558_ _06382_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__a22o_1
X_35883_ clknet_leaf_400_CLK _03997_ VGND VGND VPWR VPWR registers\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34834_ clknet_leaf_100_CLK _02948_ VGND VGND VPWR VPWR registers\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 DW[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_8
X_19768_ registers\[20\]\[39\] registers\[21\]\[39\] registers\[22\]\[39\] registers\[23\]\[39\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__mux4_1
XFILLER_231_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18719_ registers\[44\]\[10\] registers\[45\]\[10\] registers\[46\]\[10\] registers\[47\]\[10\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__mux4_1
X_34765_ clknet_leaf_148_CLK _02879_ VGND VGND VPWR VPWR registers\[25\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19699_ _06403_ _06410_ _06417_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__or4_2
X_31977_ clknet_leaf_21_CLK _00147_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21730_ registers\[56\]\[30\] registers\[57\]\[30\] registers\[58\]\[30\] registers\[59\]\[30\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__mux4_1
X_33716_ clknet_leaf_346_CLK _01830_ VGND VGND VPWR VPWR registers\[41\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30928_ registers\[10\]\[27\] _12991_ _13944_ VGND VGND VPWR VPWR _13952_ sky130_fd_sc_hd__mux2_1
X_34696_ clknet_leaf_218_CLK _02810_ VGND VGND VPWR VPWR registers\[26\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33647_ clknet_leaf_359_CLK _01761_ VGND VGND VPWR VPWR registers\[42\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_21661_ _07285_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__buf_4
X_30859_ _13915_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__clkbuf_1
X_23400_ _09854_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
X_20612_ _07292_ _07308_ _07310_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24380_ registers\[57\]\[43\] _10395_ _10389_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__mux2_1
XFILLER_51_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33578_ clknet_leaf_428_CLK _01692_ VGND VGND VPWR VPWR registers\[43\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_21592_ _07991_ _08261_ _08264_ _07995_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__a22o_1
XFILLER_123_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23331_ registers\[9\]\[58\] _09815_ _09798_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__mux2_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35317_ clknet_leaf_418_CLK _03431_ VGND VGND VPWR VPWR registers\[16\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_20543_ _07222_ _07229_ _07236_ _07243_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__or4_1
X_32529_ clknet_leaf_76_CLK _00643_ VGND VGND VPWR VPWR registers\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_37_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_37_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26050_ _10770_ registers\[45\]\[19\] _11312_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35248_ clknet_leaf_393_CLK _03362_ VGND VGND VPWR VPWR registers\[17\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_23262_ registers\[9\]\[37\] _09769_ _09754_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__mux2_1
X_20474_ _05060_ _07175_ _07176_ _05066_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__a22o_1
X_25001_ net34 VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__buf_4
X_22213_ registers\[20\]\[43\] registers\[21\]\[43\] registers\[22\]\[43\] registers\[23\]\[43\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__mux4_1
X_35179_ clknet_leaf_408_CLK _03293_ VGND VGND VPWR VPWR registers\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_23193_ registers\[9\]\[14\] _09687_ _09722_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22144_ _08766_ _08800_ _08801_ _08771_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__a22o_1
XTAP_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29740_ registers\[1\]\[40\] _13018_ _13326_ VGND VGND VPWR VPWR _13327_ sky130_fd_sc_hd__mux2_1
XTAP_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26952_ _11817_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__clkbuf_1
X_22075_ _08462_ _08732_ _08733_ _08467_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__a22o_1
XFILLER_248_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21026_ _07640_ _07713_ _07714_ _07646_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__a22o_1
X_25903_ _10758_ registers\[46\]\[13\] _11241_ VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__mux2_1
X_29671_ _13290_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__clkbuf_1
X_26883_ _11770_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_1
X_28622_ _12707_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25834_ _11208_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28553_ _12671_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__clkbuf_1
X_25765_ _11172_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
X_22977_ _09580_ registers\[62\]\[31\] _09578_ VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__mux2_1
XFILLER_215_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27504_ _12118_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__clkbuf_1
X_24716_ _10583_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28484_ _11839_ registers\[28\]\[52\] _12632_ VGND VGND VPWR VPWR _12635_ sky130_fd_sc_hd__mux2_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21928_ _08588_ _08591_ _08430_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__o21ba_1
X_25696_ registers\[48\]\[44\] _10397_ _11130_ VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27435_ _12082_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _09577_ registers\[55\]\[30\] _10547_ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__mux2_1
X_21859_ registers\[28\]\[33\] registers\[29\]\[33\] registers\[30\]\[33\] registers\[31\]\[33\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__mux4_1
XFILLER_187_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27366_ registers\[36\]\[35\] _10378_ _12040_ VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__mux2_1
X_24578_ _10509_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29105_ registers\[23\]\[17\] _12970_ _12956_ VGND VGND VPWR VPWR _12971_ sky130_fd_sc_hd__mux2_1
XFILLER_169_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26317_ _11462_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
X_23529_ _09923_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27297_ registers\[36\]\[2\] _10309_ _12007_ VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_28_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_28_CLK sky130_fd_sc_hd__clkbuf_16
X_29036_ registers\[24\]\[58\] _10426_ _12916_ VGND VGND VPWR VPWR _12925_ sky130_fd_sc_hd__mux2_1
X_17050_ _15334_ _15534_ _15535_ _15339_ VGND VGND VPWR VPWR _15536_ sky130_fd_sc_hd__a22o_1
X_26248_ _10833_ registers\[44\]\[49\] _11416_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__mux2_1
X_16001_ net68 net67 VGND VGND VPWR VPWR _14515_ sky130_fd_sc_hd__nor2b_4
XFILLER_87_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26179_ _10764_ registers\[44\]\[16\] _11383_ VGND VGND VPWR VPWR _11390_ sky130_fd_sc_hd__mux2_1
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_989 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _04722_ _04725_ _04619_ _04620_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__o211a_1
X_29938_ registers\[17\]\[6\] _12947_ _13424_ VGND VGND VPWR VPWR _13431_ sky130_fd_sc_hd__mux2_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16903_ registers\[24\]\[23\] registers\[25\]\[23\] registers\[26\]\[23\] registers\[27\]\[23\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15394_ sky130_fd_sc_hd__mux4_1
XFILLER_191_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17883_ _04548_ _04657_ _04658_ _04552_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a22o_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29869_ _13394_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31900_ _14418_ VGND VGND VPWR VPWR _14463_ sky130_fd_sc_hd__buf_4
XFILLER_152_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19622_ registers\[24\]\[35\] registers\[25\]\[35\] registers\[26\]\[35\] registers\[27\]\[35\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__mux4_1
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16834_ registers\[16\]\[21\] registers\[17\]\[21\] registers\[18\]\[21\] registers\[19\]\[21\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15327_ sky130_fd_sc_hd__mux4_1
X_32880_ clknet_leaf_368_CLK _00994_ VGND VGND VPWR VPWR registers\[54\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31831_ _09672_ registers\[49\]\[7\] _14419_ VGND VGND VPWR VPWR _14427_ sky130_fd_sc_hd__mux2_1
XFILLER_19_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19553_ registers\[4\]\[33\] registers\[5\]\[33\] registers\[6\]\[33\] registers\[7\]\[33\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__mux4_1
XFILLER_150_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16765_ _15238_ _15245_ _15252_ _15259_ VGND VGND VPWR VPWR _15260_ sky130_fd_sc_hd__or4_2
XFILLER_53_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18504_ _05240_ _05247_ _05256_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__or4_4
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34550_ clknet_leaf_313_CLK _02664_ VGND VGND VPWR VPWR registers\[28\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_234_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19484_ _06036_ _06214_ _06215_ _06039_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__a22o_1
X_31762_ _14390_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__clkbuf_1
X_16696_ registers\[32\]\[18\] registers\[33\]\[18\] registers\[34\]\[18\] registers\[35\]\[18\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15192_ sky130_fd_sc_hd__mux4_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33501_ clknet_leaf_31_CLK _01615_ VGND VGND VPWR VPWR registers\[44\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_30713_ registers\[12\]\[53\] _13046_ _13835_ VGND VGND VPWR VPWR _13839_ sky130_fd_sc_hd__mux2_1
X_18435_ _05196_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__clkbuf_1
X_34481_ clknet_leaf_385_CLK _02595_ VGND VGND VPWR VPWR registers\[2\]\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31693_ _14354_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__clkbuf_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36220_ clknet_leaf_116_CLK _00104_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dfxtp_1
X_33432_ clknet_leaf_31_CLK _01546_ VGND VGND VPWR VPWR registers\[45\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18366_ registers\[4\]\[0\] registers\[5\]\[0\] registers\[6\]\[0\] registers\[7\]\[0\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__mux4_1
X_30644_ registers\[12\]\[20\] _12976_ _13802_ VGND VGND VPWR VPWR _13803_ sky130_fd_sc_hd__mux2_1
XFILLER_226_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17317_ _15482_ _15794_ _15795_ _15485_ VGND VGND VPWR VPWR _15796_ sky130_fd_sc_hd__a22o_1
X_36151_ clknet_leaf_335_CLK _04265_ VGND VGND VPWR VPWR registers\[49\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_33363_ clknet_leaf_125_CLK _01477_ VGND VGND VPWR VPWR registers\[46\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_30575_ _13766_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__clkbuf_1
X_18297_ _05059_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__buf_4
XFILLER_30_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_19_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_222_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35102_ clknet_leaf_487_CLK _03216_ VGND VGND VPWR VPWR registers\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32314_ clknet_leaf_185_CLK _00428_ VGND VGND VPWR VPWR registers\[19\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_17248_ registers\[0\]\[33\] registers\[1\]\[33\] registers\[2\]\[33\] registers\[3\]\[33\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15729_ sky130_fd_sc_hd__mux4_1
X_36082_ clknet_leaf_363_CLK _04196_ VGND VGND VPWR VPWR registers\[59\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_33294_ clknet_leaf_130_CLK _01408_ VGND VGND VPWR VPWR registers\[47\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35033_ clknet_leaf_3_CLK _03147_ VGND VGND VPWR VPWR registers\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32245_ clknet_leaf_350_CLK _00359_ VGND VGND VPWR VPWR registers\[39\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_17179_ registers\[8\]\[31\] registers\[9\]\[31\] registers\[10\]\[31\] registers\[11\]\[31\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15662_ sky130_fd_sc_hd__mux4_1
XFILLER_31_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20190_ _06722_ _06900_ _06901_ _06725_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__a22o_1
XFILLER_116_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32176_ clknet_leaf_14_CLK _00290_ VGND VGND VPWR VPWR registers\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31127_ _14056_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35935_ clknet_leaf_480_CLK _04049_ VGND VGND VPWR VPWR registers\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_31058_ _14020_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22900_ _09528_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
X_30009_ _13423_ VGND VGND VPWR VPWR _13468_ sky130_fd_sc_hd__buf_4
XFILLER_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23880_ _10088_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__buf_4
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35866_ clknet_leaf_476_CLK _03980_ VGND VGND VPWR VPWR registers\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22831_ _07276_ _09466_ _09467_ _07286_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__a22o_1
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34817_ clknet_leaf_225_CLK _02931_ VGND VGND VPWR VPWR registers\[24\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_35797_ clknet_leaf_79_CLK _03911_ VGND VGND VPWR VPWR registers\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_909 _09689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22762_ registers\[56\]\[60\] registers\[57\]\[60\] registers\[58\]\[60\] registers\[59\]\[60\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__mux4_1
X_25550_ registers\[4\]\[40\] _10388_ _11056_ VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__mux2_1
X_34748_ clknet_leaf_188_CLK _02862_ VGND VGND VPWR VPWR registers\[25\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21713_ _08075_ _08381_ _08382_ _08078_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__a22o_1
X_24501_ _10469_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
X_25481_ _11020_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22693_ _09313_ _09320_ _09327_ _09334_ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__or4_4
XFILLER_129_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34679_ clknet_leaf_311_CLK _02793_ VGND VGND VPWR VPWR registers\[26\]\[41\] sky130_fd_sc_hd__dfxtp_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27220_ _11935_ VGND VGND VPWR VPWR _11969_ sky130_fd_sc_hd__buf_4
XFILLER_205_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24432_ registers\[57\]\[60\] _10430_ net283 VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__mux2_1
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21644_ _08080_ _08314_ _08315_ _08085_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__a22o_1
XFILLER_240_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27151_ _11932_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24363_ net32 VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__buf_4
XFILLER_21_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_40 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ _08245_ _08248_ _08087_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__o21ba_1
XFILLER_201_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_51 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23314_ registers\[9\]\[53\] _09804_ _09798_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__mux2_1
X_26102_ _11349_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_62 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20526_ registers\[52\]\[62\] registers\[53\]\[62\] registers\[54\]\[62\] registers\[55\]\[62\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__mux4_1
XANTENNA_73 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27082_ _11896_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_84 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24294_ _10337_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_95 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26033_ _11313_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
X_23245_ registers\[9\]\[32\] _09758_ _09754_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__mux2_1
X_20457_ _06912_ _07158_ _07159_ _06917_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__a22o_1
XFILLER_10_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23176_ registers\[39\]\[22\] _09717_ _09700_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__mux2_1
X_20388_ _06868_ _07092_ _07093_ _06871_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__a22o_1
XFILLER_175_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22127_ _08669_ _08783_ _08784_ _08675_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__a22o_1
XTAP_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1308 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27984_ _11744_ registers\[31\]\[7\] _12364_ VGND VGND VPWR VPWR _12372_ sky130_fd_sc_hd__mux2_1
XANTENNA_1319 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput180 net180 VGND VGND VPWR VPWR D2[33] sky130_fd_sc_hd__buf_2
XFILLER_216_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput191 net191 VGND VGND VPWR VPWR D2[43] sky130_fd_sc_hd__buf_2
XTAP_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29723_ registers\[1\]\[32\] _13002_ _13315_ VGND VGND VPWR VPWR _13318_ sky130_fd_sc_hd__mux2_1
XTAP_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26935_ _11805_ registers\[3\]\[36\] _11793_ VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__mux2_1
X_22058_ registers\[0\]\[39\] registers\[1\]\[39\] registers\[2\]\[39\] registers\[3\]\[39\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__mux4_1
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21009_ registers\[20\]\[9\] registers\[21\]\[9\] registers\[22\]\[9\] registers\[23\]\[9\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__mux4_1
X_29654_ _09707_ _11008_ VGND VGND VPWR VPWR _13281_ sky130_fd_sc_hd__nor2_8
XTAP_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26866_ net6 VGND VGND VPWR VPWR _11759_ sky130_fd_sc_hd__buf_4
XTAP_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28605_ _12698_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25817_ _11199_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
X_29585_ _13245_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26797_ registers\[40\]\[52\] _10414_ _11713_ VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__mux2_1
XFILLER_56_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28536_ _12662_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__clkbuf_1
X_16550_ registers\[24\]\[13\] registers\[25\]\[13\] registers\[26\]\[13\] registers\[27\]\[13\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _15051_ sky130_fd_sc_hd__mux4_1
X_25748_ _11163_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28467_ _11822_ registers\[28\]\[44\] _12621_ VGND VGND VPWR VPWR _12626_ sky130_fd_sc_hd__mux2_1
X_16481_ registers\[16\]\[11\] registers\[17\]\[11\] registers\[18\]\[11\] registers\[19\]\[11\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14984_ sky130_fd_sc_hd__mux4_1
XFILLER_204_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25679_ registers\[48\]\[36\] _10380_ _11119_ VGND VGND VPWR VPWR _11126_ sky130_fd_sc_hd__mux2_1
XFILLER_204_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18220_ _14540_ _04983_ _04984_ _14551_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a22o_1
XFILLER_70_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27418_ registers\[36\]\[60\] _10430_ _12006_ VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28398_ _11753_ registers\[28\]\[11\] _12588_ VGND VGND VPWR VPWR _12590_ sky130_fd_sc_hd__mux2_1
XFILLER_70_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18151_ _04637_ _04917_ _04918_ _04642_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__a22o_1
X_27349_ registers\[36\]\[27\] _10361_ _12029_ VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__mux2_1
XFILLER_223_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17102_ _15549_ _15585_ _15586_ _15553_ VGND VGND VPWR VPWR _15587_ sky130_fd_sc_hd__a22o_1
XFILLER_89_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18082_ registers\[12\]\[57\] registers\[13\]\[57\] registers\[14\]\[57\] registers\[15\]\[57\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__mux4_1
X_30360_ _13653_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29019_ _12860_ VGND VGND VPWR VPWR _12916_ sky130_fd_sc_hd__buf_4
XFILLER_221_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17033_ registers\[0\]\[27\] registers\[1\]\[27\] registers\[2\]\[27\] registers\[3\]\[27\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15520_ sky130_fd_sc_hd__mux4_1
X_30291_ _13616_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32030_ clknet_leaf_50_CLK _00208_ VGND VGND VPWR VPWR registers\[62\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _05693_ _05728_ _05729_ _05696_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__a22o_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17935_ _04637_ _04708_ _04709_ _04642_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a22o_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33981_ clknet_leaf_268_CLK _02095_ VGND VGND VPWR VPWR registers\[37\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35720_ clknet_leaf_154_CLK _03834_ VGND VGND VPWR VPWR registers\[10\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32932_ clknet_leaf_442_CLK _01046_ VGND VGND VPWR VPWR registers\[53\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17866_ _04637_ _04638_ _04641_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_8_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_8_CLK sky130_fd_sc_hd__clkbuf_16
X_19605_ _06329_ _06332_ _06161_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__o21ba_1
X_16817_ _14998_ _15308_ _15309_ _15001_ VGND VGND VPWR VPWR _15310_ sky130_fd_sc_hd__a22o_1
X_35651_ clknet_leaf_243_CLK _03765_ VGND VGND VPWR VPWR registers\[11\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32863_ clknet_leaf_45_CLK _00977_ VGND VGND VPWR VPWR registers\[54\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17797_ registers\[32\]\[49\] registers\[33\]\[49\] registers\[34\]\[49\] registers\[35\]\[49\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__mux4_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31814_ _14417_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__clkbuf_1
X_19536_ registers\[44\]\[33\] registers\[45\]\[33\] registers\[46\]\[33\] registers\[47\]\[33\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux4_1
X_34602_ clknet_leaf_407_CLK _02716_ VGND VGND VPWR VPWR registers\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_35582_ clknet_leaf_297_CLK _03696_ VGND VGND VPWR VPWR registers\[12\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16748_ registers\[52\]\[19\] registers\[53\]\[19\] registers\[54\]\[19\] registers\[55\]\[19\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15243_ sky130_fd_sc_hd__mux4_1
XFILLER_228_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32794_ clknet_leaf_67_CLK _00908_ VGND VGND VPWR VPWR registers\[55\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_34533_ clknet_leaf_456_CLK _02647_ VGND VGND VPWR VPWR registers\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31745_ registers\[59\]\[30\] net24 _14381_ VGND VGND VPWR VPWR _14382_ sky130_fd_sc_hd__mux2_1
X_19467_ _05883_ _06197_ _06198_ _05888_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__a22o_1
X_16679_ registers\[8\]\[17\] registers\[9\]\[17\] registers\[10\]\[17\] registers\[11\]\[17\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15176_ sky130_fd_sc_hd__mux4_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18418_ _05089_ _05178_ _05179_ _05100_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__a22o_1
X_34464_ clknet_leaf_487_CLK _02578_ VGND VGND VPWR VPWR registers\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31676_ registers\[63\]\[62\] net59 _14276_ VGND VGND VPWR VPWR _14345_ sky130_fd_sc_hd__mux2_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19398_ registers\[48\]\[29\] registers\[49\]\[29\] registers\[50\]\[29\] registers\[51\]\[29\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__mux4_1
XFILLER_194_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33415_ clknet_leaf_251_CLK _01529_ VGND VGND VPWR VPWR registers\[46\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_36203_ clknet_leaf_22_CLK _00085_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dfxtp_2
X_18349_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__buf_6
X_30627_ registers\[12\]\[12\] _12960_ _13791_ VGND VGND VPWR VPWR _13794_ sky130_fd_sc_hd__mux2_1
X_34395_ clknet_leaf_1_CLK _02509_ VGND VGND VPWR VPWR registers\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36134_ clknet_leaf_434_CLK _04248_ VGND VGND VPWR VPWR registers\[49\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_33346_ clknet_leaf_256_CLK _01460_ VGND VGND VPWR VPWR registers\[47\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_21360_ _07732_ _08038_ _08039_ _07735_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__a22o_1
XFILLER_174_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30558_ _13757_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20311_ _07015_ _07018_ _06847_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__o21ba_1
XFILLER_200_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36065_ clknet_leaf_43_CLK _04179_ VGND VGND VPWR VPWR registers\[59\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_33277_ clknet_leaf_283_CLK _01391_ VGND VGND VPWR VPWR registers\[48\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_21291_ _07737_ _07971_ _07972_ _07742_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__a22o_1
Xinput60 DW[63] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_16
Xinput71 R2[0] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30489_ _13721_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__clkbuf_1
Xinput82 R3[5] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
X_35016_ clknet_leaf_208_CLK _03130_ VGND VGND VPWR VPWR registers\[21\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_23030_ _09616_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
X_32228_ clknet_leaf_154_CLK _00342_ VGND VGND VPWR VPWR registers\[9\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_20242_ registers\[44\]\[53\] registers\[45\]\[53\] registers\[46\]\[53\] registers\[47\]\[53\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__mux4_1
XFILLER_200_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20173_ _06569_ _06883_ _06884_ _06574_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__a22o_1
XFILLER_153_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32159_ clknet_leaf_40_CLK _00273_ VGND VGND VPWR VPWR registers\[39\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24981_ _09640_ registers\[53\]\[60\] _10657_ VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26720_ _11675_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35918_ clknet_leaf_138_CLK _04032_ VGND VGND VPWR VPWR registers\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ _10138_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26651_ _11638_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__clkbuf_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35849_ clknet_leaf_155_CLK _03963_ VGND VGND VPWR VPWR registers\[8\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_23863_ _10102_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25602_ _11082_ _11084_ VGND VGND VPWR VPWR _11085_ sky130_fd_sc_hd__nor2_8
XANTENNA_706 _07287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22814_ _09451_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
X_29370_ _09813_ registers\[22\]\[57\] _13124_ VGND VGND VPWR VPWR _13132_ sky130_fd_sc_hd__mux2_1
XANTENNA_717 _07312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_728 _07349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26582_ _11602_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_739 _07359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23794_ _10065_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28321_ registers\[2\]\[39\] _10386_ _12539_ VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__mux2_1
X_25533_ registers\[4\]\[32\] _10372_ _11045_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22745_ _09381_ _09384_ _09102_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__o21ba_1
XFILLER_207_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28252_ registers\[2\]\[6\] _10317_ _12506_ VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__mux2_1
XFILLER_13_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25464_ _11008_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__nor2_8
XFILLER_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22676_ registers\[52\]\[57\] registers\[53\]\[57\] registers\[54\]\[57\] registers\[55\]\[57\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27203_ _11960_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__clkbuf_1
X_24415_ _10419_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21627_ _07983_ _08297_ _08298_ _07989_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__a22o_1
X_28183_ _12476_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__clkbuf_1
X_25395_ _10973_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27134_ _11841_ registers\[38\]\[53\] _11920_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__mux2_1
X_24346_ registers\[57\]\[32\] _10372_ _10368_ VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__mux2_1
X_21558_ _07991_ _08230_ _08231_ _07995_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__a22o_1
XFILLER_153_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20509_ registers\[28\]\[61\] registers\[29\]\[61\] registers\[30\]\[61\] registers\[31\]\[61\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__mux4_1
X_24277_ net283 VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__clkbuf_8
X_27065_ _11771_ registers\[38\]\[20\] _11887_ VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__mux2_1
X_21489_ _07983_ _08163_ _08164_ _07989_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26016_ _11304_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
XTAP_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23228_ net20 VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23159_ _09705_ _09707_ VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__nor2_8
XTAP_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1105 _14553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1116 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1127 _14597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1138 _14613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15981_ net66 VGND VGND VPWR VPWR _14495_ sky130_fd_sc_hd__clkbuf_16
XTAP_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27967_ _12362_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1149 _15676_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _04471_ _04480_ _04491_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__or4_4
X_29706_ registers\[1\]\[24\] _12985_ _13304_ VGND VGND VPWR VPWR _13309_ sky130_fd_sc_hd__mux2_1
XTAP_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26918_ _11794_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27898_ registers\[32\]\[30\] _10367_ _12326_ VGND VGND VPWR VPWR _12327_ sky130_fd_sc_hd__mux2_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29637_ _13272_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__clkbuf_1
XTAP_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _04433_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkbuf_4
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26849_ _11747_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _14855_ _15099_ _15100_ _14861_ VGND VGND VPWR VPWR _15101_ sky130_fd_sc_hd__a22o_1
X_17582_ _04294_ _04365_ _04366_ _04299_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__a22o_1
X_29568_ _13236_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19321_ _05122_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__buf_4
XFILLER_216_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28519_ _12653_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__clkbuf_1
X_16533_ _15030_ _15033_ _14926_ VGND VGND VPWR VPWR _15034_ sky130_fd_sc_hd__o21ba_1
X_29499_ _09806_ registers\[21\]\[54\] _13195_ VGND VGND VPWR VPWR _13200_ sky130_fd_sc_hd__mux2_1
XFILLER_56_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31530_ _14268_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__clkbuf_1
X_19252_ _05986_ _05989_ _05818_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__o21ba_1
XFILLER_232_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16464_ _14655_ _14965_ _14966_ _14658_ VGND VGND VPWR VPWR _14967_ sky130_fd_sc_hd__a22o_1
XFILLER_177_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18203_ registers\[4\]\[61\] registers\[5\]\[61\] registers\[6\]\[61\] registers\[7\]\[61\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__mux4_1
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19183_ registers\[44\]\[23\] registers\[45\]\[23\] registers\[46\]\[23\] registers\[47\]\[23\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__mux4_1
X_31461_ _14232_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__clkbuf_1
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16395_ registers\[52\]\[9\] registers\[53\]\[9\] registers\[54\]\[9\] registers\[55\]\[9\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14900_ sky130_fd_sc_hd__mux4_1
XFILLER_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33200_ clknet_leaf_373_CLK _01314_ VGND VGND VPWR VPWR registers\[4\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_18134_ _14587_ _04900_ _04901_ _14597_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__a22o_1
X_30412_ _13680_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__clkbuf_1
X_34180_ clknet_leaf_246_CLK _02294_ VGND VGND VPWR VPWR registers\[34\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31392_ registers\[7\]\[55\] net51 _14190_ VGND VGND VPWR VPWR _14196_ sky130_fd_sc_hd__mux2_1
XFILLER_172_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33131_ clknet_leaf_425_CLK _01245_ VGND VGND VPWR VPWR registers\[50\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_18065_ registers\[40\]\[57\] registers\[41\]\[57\] registers\[42\]\[57\] registers\[43\]\[57\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__mux4_1
X_30343_ _13644_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17016_ registers\[40\]\[27\] registers\[41\]\[27\] registers\[42\]\[27\] registers\[43\]\[27\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15503_ sky130_fd_sc_hd__mux4_1
XFILLER_172_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33062_ clknet_leaf_439_CLK _01176_ VGND VGND VPWR VPWR registers\[51\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_30274_ _13607_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32013_ clknet_leaf_92_CLK _00187_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18967_ _05120_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__buf_4
XFILLER_112_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1650 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1090 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1661 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1672 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17918_ registers\[52\]\[52\] registers\[53\]\[52\] registers\[54\]\[52\] registers\[55\]\[52\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__mux4_1
XFILLER_227_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1683 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33964_ clknet_leaf_325_CLK _02078_ VGND VGND VPWR VPWR registers\[37\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_18898_ _05547_ _05644_ _05645_ _05550_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__a22o_1
XANTENNA_1694 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35703_ clknet_leaf_318_CLK _03817_ VGND VGND VPWR VPWR registers\[10\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_17849_ _04481_ _04622_ _04625_ _04484_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__a22o_1
X_32915_ clknet_leaf_182_CLK _01029_ VGND VGND VPWR VPWR registers\[53\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_33895_ clknet_leaf_434_CLK _02009_ VGND VGND VPWR VPWR registers\[38\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20860_ registers\[4\]\[5\] registers\[5\]\[5\] registers\[6\]\[5\] registers\[7\]\[5\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__mux4_1
X_32846_ clknet_leaf_180_CLK _00960_ VGND VGND VPWR VPWR registers\[54\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_35634_ clknet_leaf_381_CLK _03748_ VGND VGND VPWR VPWR registers\[11\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19519_ registers\[4\]\[32\] registers\[5\]\[32\] registers\[6\]\[32\] registers\[7\]\[32\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__mux4_1
XFILLER_74_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32777_ clknet_leaf_210_CLK _00891_ VGND VGND VPWR VPWR registers\[56\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20791_ _07356_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__buf_6
X_35565_ clknet_leaf_392_CLK _03679_ VGND VGND VPWR VPWR registers\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_250_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_250_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22530_ _09104_ _09175_ _09176_ _09107_ VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__a22o_1
XFILLER_168_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34516_ clknet_leaf_94_CLK _02630_ VGND VGND VPWR VPWR registers\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31728_ registers\[59\]\[22\] net15 _14370_ VGND VGND VPWR VPWR _14373_ sky130_fd_sc_hd__mux2_1
X_35496_ clknet_leaf_398_CLK _03610_ VGND VGND VPWR VPWR registers\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22461_ registers\[28\]\[50\] registers\[29\]\[50\] registers\[30\]\[50\] registers\[31\]\[50\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__mux4_1
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34447_ clknet_leaf_110_CLK _02561_ VGND VGND VPWR VPWR registers\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_31659_ _14336_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24200_ _10280_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
X_21412_ registers\[40\]\[21\] registers\[41\]\[21\] registers\[42\]\[21\] registers\[43\]\[21\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__mux4_1
X_25180_ net58 VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__buf_2
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34378_ clknet_leaf_166_CLK _02492_ VGND VGND VPWR VPWR registers\[31\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_22392_ _09011_ _09026_ _09035_ _09042_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__or4_4
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24131_ _10232_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__buf_6
X_36117_ clknet_leaf_70_CLK _04231_ VGND VGND VPWR VPWR registers\[49\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_33329_ clknet_leaf_361_CLK _01443_ VGND VGND VPWR VPWR registers\[47\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_21343_ _08019_ _08022_ _07711_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__o21ba_1
X_24062_ _10207_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__clkbuf_1
X_36048_ clknet_leaf_73_CLK _04162_ VGND VGND VPWR VPWR registers\[59\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_21274_ _07640_ _07954_ _07955_ _07646_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__a22o_1
XFILLER_150_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23013_ net38 VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_239_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20225_ registers\[4\]\[52\] registers\[5\]\[52\] registers\[6\]\[52\] registers\[7\]\[52\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__mux4_1
X_28870_ _11820_ registers\[25\]\[43\] _12834_ VGND VGND VPWR VPWR _12838_ sky130_fd_sc_hd__mux2_1
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27821_ registers\[33\]\[58\] _10426_ _12277_ VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__mux2_1
XFILLER_133_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20156_ registers\[24\]\[50\] registers\[25\]\[50\] registers\[26\]\[50\] registers\[27\]\[50\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__mux4_1
XFILLER_131_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27752_ registers\[33\]\[25\] _10357_ _12244_ VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__mux2_1
XFILLER_246_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24964_ _10715_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__clkbuf_1
X_20087_ _06525_ _06800_ _06801_ _06528_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__a22o_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26703_ _11666_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_1
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _10129_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
X_27683_ _12213_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_218_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24895_ _09554_ registers\[53\]\[19\] _10669_ VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__mux2_1
XFILLER_73_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29422_ _13159_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__clkbuf_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26634_ _11629_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_503 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23846_ _10093_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__clkbuf_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_514 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_525 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29353_ _09795_ registers\[22\]\[49\] _13113_ VGND VGND VPWR VPWR _13123_ sky130_fd_sc_hd__mux2_1
XANTENNA_547 _04345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26565_ _11593_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_558 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _07440_ _07677_ _07678_ _07443_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__a22o_1
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23777_ _10056_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_569 _04834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_241_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_241_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28304_ _12540_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__clkbuf_1
X_25516_ registers\[4\]\[24\] _10355_ _11034_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__mux2_1
X_22728_ registers\[44\]\[59\] registers\[45\]\[59\] registers\[46\]\[59\] registers\[47\]\[59\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__mux4_1
X_29284_ _09691_ registers\[22\]\[16\] _13080_ VGND VGND VPWR VPWR _13087_ sky130_fd_sc_hd__mux2_1
X_26496_ _11556_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
X_28235_ _12503_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25447_ _11000_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22659_ registers\[28\]\[56\] registers\[29\]\[56\] registers\[30\]\[56\] registers\[31\]\[56\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__mux4_1
XFILLER_16_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16180_ _14687_ _14690_ _14525_ VGND VGND VPWR VPWR _14691_ sky130_fd_sc_hd__o21ba_1
X_28166_ _12467_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25378_ _10964_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27117_ _11824_ registers\[38\]\[45\] _11909_ VGND VGND VPWR VPWR _11915_ sky130_fd_sc_hd__mux2_1
X_24329_ net20 VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__buf_4
X_28097_ _11857_ registers\[31\]\[61\] _12363_ VGND VGND VPWR VPWR _12431_ sky130_fd_sc_hd__mux2_1
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27048_ _11755_ registers\[38\]\[12\] _11876_ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__mux2_1
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19870_ _06374_ _06589_ _06590_ _06377_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__a22o_1
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18821_ registers\[28\]\[12\] registers\[29\]\[12\] registers\[30\]\[12\] registers\[31\]\[12\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__mux4_1
XTAP_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28999_ registers\[24\]\[40\] _10388_ _12905_ VGND VGND VPWR VPWR _12906_ sky130_fd_sc_hd__mux2_1
XTAP_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18752_ registers\[20\]\[10\] registers\[21\]\[10\] registers\[22\]\[10\] registers\[23\]\[10\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__mux4_1
XTAP_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17703_ _14567_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__buf_4
XFILLER_248_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18683_ _05067_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__buf_6
X_30961_ _13969_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32700_ clknet_leaf_284_CLK _00814_ VGND VGND VPWR VPWR registers\[57\]\[46\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_480_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_480_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ registers\[8\]\[44\] registers\[9\]\[44\] registers\[10\]\[44\] registers\[11\]\[44\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__mux4_1
X_33680_ clknet_leaf_129_CLK _01794_ VGND VGND VPWR VPWR registers\[41\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30892_ _13921_ VGND VGND VPWR VPWR _13933_ sky130_fd_sc_hd__buf_4
X_32631_ clknet_leaf_328_CLK _00745_ VGND VGND VPWR VPWR registers\[58\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17565_ registers\[52\]\[42\] registers\[53\]\[42\] registers\[54\]\[42\] registers\[55\]\[42\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_232_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_232_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19304_ _06035_ _06040_ _05837_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__o21ba_1
XFILLER_90_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35350_ clknet_leaf_82_CLK _03464_ VGND VGND VPWR VPWR registers\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_16516_ registers\[24\]\[12\] registers\[25\]\[12\] registers\[26\]\[12\] registers\[27\]\[12\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _15018_ sky130_fd_sc_hd__mux4_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32562_ clknet_leaf_379_CLK _00676_ VGND VGND VPWR VPWR registers\[5\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17496_ _15825_ _15966_ _15969_ _15828_ VGND VGND VPWR VPWR _15970_ sky130_fd_sc_hd__a22o_1
X_31513_ _14259_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__clkbuf_1
X_34301_ clknet_leaf_277_CLK _02415_ VGND VGND VPWR VPWR registers\[32\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19235_ _05111_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__buf_6
X_35281_ clknet_leaf_106_CLK _03395_ VGND VGND VPWR VPWR registers\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16447_ _14947_ _14948_ _14949_ _14950_ VGND VGND VPWR VPWR _14951_ sky130_fd_sc_hd__a22o_1
X_32493_ clknet_leaf_374_CLK _00607_ VGND VGND VPWR VPWR registers\[60\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34232_ clknet_leaf_338_CLK _02346_ VGND VGND VPWR VPWR registers\[33\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_19166_ registers\[4\]\[22\] registers\[5\]\[22\] registers\[6\]\[22\] registers\[7\]\[22\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__mux4_1
X_31444_ _14223_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16378_ _14601_ _14882_ _14883_ _14611_ VGND VGND VPWR VPWR _14884_ sky130_fd_sc_hd__a22o_1
XFILLER_129_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18117_ registers\[16\]\[58\] registers\[17\]\[58\] registers\[18\]\[58\] registers\[19\]\[58\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__mux4_1
XFILLER_160_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34163_ clknet_leaf_349_CLK _02277_ VGND VGND VPWR VPWR registers\[34\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31375_ registers\[7\]\[47\] net42 _14179_ VGND VGND VPWR VPWR _14187_ sky130_fd_sc_hd__mux2_1
X_19097_ registers\[24\]\[20\] registers\[25\]\[20\] registers\[26\]\[20\] registers\[27\]\[20\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33114_ clknet_leaf_84_CLK _01228_ VGND VGND VPWR VPWR registers\[50\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_30326_ _13634_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__clkbuf_1
X_18048_ _04815_ _04818_ _04619_ _04620_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__o211a_1
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34094_ clknet_leaf_355_CLK _02208_ VGND VGND VPWR VPWR registers\[35\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_299_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_299_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33045_ clknet_leaf_69_CLK _01159_ VGND VGND VPWR VPWR registers\[51\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_30257_ _13598_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20010_ _06721_ _06726_ _06523_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__o21ba_1
XFILLER_28_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30188_ registers\[16\]\[61\] _13062_ _13494_ VGND VGND VPWR VPWR _13562_ sky130_fd_sc_hd__mux2_1
XFILLER_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19999_ _06710_ _06715_ _06512_ _06513_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__o211a_1
XFILLER_80_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34996_ clknet_leaf_414_CLK _03110_ VGND VGND VPWR VPWR registers\[21\]\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1480 _05654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1491 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21961_ registers\[16\]\[36\] registers\[17\]\[36\] registers\[18\]\[36\] registers\[19\]\[36\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__mux4_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33947_ clknet_leaf_24_CLK _02061_ VGND VGND VPWR VPWR registers\[37\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23700_ _09654_ _09941_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__nor2_8
Xclkbuf_leaf_471_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_471_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20912_ _07433_ _07602_ _07603_ _07438_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__a22o_1
X_24680_ _09611_ registers\[55\]\[46\] _10558_ VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__mux2_1
X_21892_ _08418_ _08555_ _08556_ _08421_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__a22o_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33878_ clknet_leaf_117_CLK _01992_ VGND VGND VPWR VPWR registers\[38\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ registers\[44\]\[5\] registers\[45\]\[5\] registers\[46\]\[5\] registers\[47\]\[5\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__mux4_1
X_23631_ _09978_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
X_35617_ clknet_leaf_485_CLK _03731_ VGND VGND VPWR VPWR registers\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32829_ clknet_leaf_289_CLK _00943_ VGND VGND VPWR VPWR registers\[55\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_223_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_223_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26350_ _10800_ registers\[43\]\[33\] _11476_ VGND VGND VPWR VPWR _11480_ sky130_fd_sc_hd__mux2_1
X_20774_ registers\[40\]\[3\] registers\[41\]\[3\] registers\[42\]\[3\] registers\[43\]\[3\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__mux4_1
X_23562_ net84 net85 VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__nand2b_4
XFILLER_223_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35548_ clknet_leaf_477_CLK _03662_ VGND VGND VPWR VPWR registers\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25301_ _10923_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22513_ _09154_ _09159_ _09083_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26281_ _10728_ registers\[43\]\[0\] _11443_ VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__mux2_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23493_ _09580_ registers\[19\]\[31\] _09903_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__mux2_1
XFILLER_196_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35479_ clknet_leaf_82_CLK _03593_ VGND VGND VPWR VPWR registers\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28020_ _11780_ registers\[31\]\[24\] _12386_ VGND VGND VPWR VPWR _12391_ sky130_fd_sc_hd__mux2_1
XFILLER_91_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22444_ _09087_ _09090_ _09091_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__o211a_1
X_25232_ _10864_ VGND VGND VPWR VPWR _10887_ sky130_fd_sc_hd__buf_4
XFILLER_176_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25163_ _10846_ registers\[52\]\[55\] _10836_ VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__mux2_1
X_22375_ _09019_ _09025_ _08748_ _08749_ VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__o211a_1
XFILLER_163_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24114_ _10235_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__clkbuf_1
X_21326_ registers\[24\]\[18\] registers\[25\]\[18\] registers\[26\]\[18\] registers\[27\]\[18\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__mux4_1
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25094_ net27 VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__clkbuf_4
X_29971_ _13448_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28922_ _12865_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24045_ _10198_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__clkbuf_1
X_21257_ registers\[28\]\[16\] registers\[29\]\[16\] registers\[30\]\[16\] registers\[31\]\[16\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__mux4_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20208_ _05088_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__buf_4
XFILLER_137_1364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28853_ _11803_ registers\[25\]\[35\] _12823_ VGND VGND VPWR VPWR _12829_ sky130_fd_sc_hd__mux2_1
XFILLER_85_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21188_ registers\[20\]\[14\] registers\[21\]\[14\] registers\[22\]\[14\] registers\[23\]\[14\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27804_ _12221_ VGND VGND VPWR VPWR _12277_ sky130_fd_sc_hd__buf_4
X_20139_ registers\[60\]\[50\] registers\[61\]\[50\] registers\[62\]\[50\] registers\[63\]\[50\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__mux4_1
XFILLER_38_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28784_ _11734_ registers\[25\]\[2\] _12790_ VGND VGND VPWR VPWR _12793_ sky130_fd_sc_hd__mux2_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25996_ _11293_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27735_ registers\[33\]\[17\] _10340_ _12233_ VGND VGND VPWR VPWR _12241_ sky130_fd_sc_hd__mux2_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24947_ _10706_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_462_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_462_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27666_ _12204_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__clkbuf_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24878_ _10670_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_300 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_311 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29405_ _13150_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_322 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_333 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26617_ _10796_ registers\[41\]\[31\] _11619_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__mux2_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23829_ _10083_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27597_ _12168_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__clkbuf_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_355 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_214_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_214_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_366 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_377 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29336_ _13114_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__clkbuf_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17350_ _14567_ VGND VGND VPWR VPWR _15828_ sky130_fd_sc_hd__buf_4
XANTENNA_388 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26548_ _11583_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_1365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_399 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _14594_ VGND VGND VPWR VPWR _14809_ sky130_fd_sc_hd__buf_4
XFILLER_109_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29267_ _09674_ registers\[22\]\[8\] _13069_ VGND VGND VPWR VPWR _13078_ sky130_fd_sc_hd__mux2_1
X_17281_ registers\[8\]\[34\] registers\[9\]\[34\] registers\[10\]\[34\] registers\[11\]\[34\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15761_ sky130_fd_sc_hd__mux4_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26479_ _10793_ registers\[42\]\[30\] _11547_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__mux2_1
XFILLER_186_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19020_ registers\[12\]\[18\] registers\[13\]\[18\] registers\[14\]\[18\] registers\[15\]\[18\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__mux4_1
X_28218_ _11843_ registers\[30\]\[54\] _12490_ VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__mux2_1
X_16232_ registers\[16\]\[4\] registers\[17\]\[4\] registers\[18\]\[4\] registers\[19\]\[4\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14742_ sky130_fd_sc_hd__mux4_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29198_ registers\[23\]\[47\] _13033_ _13019_ VGND VGND VPWR VPWR _13034_ sky130_fd_sc_hd__mux2_1
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ registers\[24\]\[2\] registers\[25\]\[2\] registers\[26\]\[2\] registers\[27\]\[2\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _14675_ sky130_fd_sc_hd__mux4_1
X_28149_ _11774_ registers\[30\]\[21\] _12457_ VGND VGND VPWR VPWR _12459_ sky130_fd_sc_hd__mux2_1
XFILLER_166_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31160_ registers\[8\]\[9\] net64 _14064_ VGND VGND VPWR VPWR _14074_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16094_ _14607_ VGND VGND VPWR VPWR _14608_ sky130_fd_sc_hd__buf_4
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30111_ registers\[16\]\[24\] _12985_ _13517_ VGND VGND VPWR VPWR _13522_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19922_ registers\[36\]\[44\] registers\[37\]\[44\] registers\[38\]\[44\] registers\[39\]\[44\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__mux4_1
XFILLER_79_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31091_ registers\[0\]\[40\] _13018_ _14037_ VGND VGND VPWR VPWR _14038_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30042_ _13485_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__clkbuf_1
X_19853_ _05049_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18804_ _05404_ _05553_ _05554_ _05410_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__a22o_1
XFILLER_228_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34850_ clknet_leaf_473_CLK _02964_ VGND VGND VPWR VPWR registers\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_16996_ registers\[0\]\[26\] registers\[1\]\[26\] registers\[2\]\[26\] registers\[3\]\[26\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15484_ sky130_fd_sc_hd__mux4_1
X_19784_ registers\[48\]\[40\] registers\[49\]\[40\] registers\[50\]\[40\] registers\[51\]\[40\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__mux4_1
X_33801_ clknet_leaf_245_CLK _01915_ VGND VGND VPWR VPWR registers\[40\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18735_ _05113_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34781_ clknet_leaf_8_CLK _02895_ VGND VGND VPWR VPWR registers\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_31993_ clknet_leaf_23_CLK _00165_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
XFILLER_95_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_453_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_453_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33732_ clknet_leaf_250_CLK _01846_ VGND VGND VPWR VPWR registers\[41\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_18666_ _05345_ _05419_ _05420_ _05348_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a22o_1
X_30944_ _13960_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__clkbuf_1
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17617_ _04400_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_4
X_30875_ _13924_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__clkbuf_1
X_33663_ clknet_leaf_272_CLK _01777_ VGND VGND VPWR VPWR registers\[42\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_18597_ _05350_ _05351_ _05352_ _05353_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_205_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_205_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35402_ clknet_leaf_150_CLK _03516_ VGND VGND VPWR VPWR registers\[15\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17548_ _14527_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__clkbuf_4
X_32614_ clknet_leaf_438_CLK _00728_ VGND VGND VPWR VPWR registers\[58\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33594_ clknet_leaf_280_CLK _01708_ VGND VGND VPWR VPWR registers\[43\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35333_ clknet_leaf_219_CLK _03447_ VGND VGND VPWR VPWR registers\[16\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32545_ clknet_leaf_470_CLK _00659_ VGND VGND VPWR VPWR registers\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_17479_ registers\[36\]\[40\] registers\[37\]\[40\] registers\[38\]\[40\] registers\[39\]\[40\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _15953_ sky130_fd_sc_hd__mux4_1
XFILLER_221_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19218_ _05953_ _05956_ _05818_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__o21ba_1
X_35264_ clknet_leaf_222_CLK _03378_ VGND VGND VPWR VPWR registers\[17\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_20490_ _06919_ _07190_ _07191_ _06922_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__a22o_1
X_32476_ clknet_leaf_53_CLK _00590_ VGND VGND VPWR VPWR registers\[60\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31427_ _14214_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__clkbuf_1
X_19149_ _05088_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__clkbuf_4
X_34215_ clknet_leaf_431_CLK _02329_ VGND VGND VPWR VPWR registers\[33\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_35195_ clknet_leaf_185_CLK _03309_ VGND VGND VPWR VPWR registers\[18\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22160_ _08811_ _08816_ _08740_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__o21ba_1
X_34146_ clknet_leaf_49_CLK _02260_ VGND VGND VPWR VPWR registers\[34\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31358_ registers\[7\]\[39\] net33 _14168_ VGND VGND VPWR VPWR _14178_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21111_ _07581_ _07796_ _07797_ _07584_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__a22o_1
X_30309_ registers\[15\]\[54\] _13048_ _13621_ VGND VGND VPWR VPWR _13626_ sky130_fd_sc_hd__mux2_1
XFILLER_59_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34077_ clknet_leaf_22_CLK _02191_ VGND VGND VPWR VPWR registers\[35\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_22091_ _08744_ _08747_ _08748_ _08749_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__o211a_1
XTAP_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31289_ registers\[7\]\[6\] net61 _14135_ VGND VGND VPWR VPWR _14142_ sky130_fd_sc_hd__mux2_1
X_33028_ clknet_leaf_259_CLK _01142_ VGND VGND VPWR VPWR registers\[52\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21042_ _07726_ _07729_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25850_ _10840_ registers\[47\]\[52\] _11214_ VGND VGND VPWR VPWR _11217_ sky130_fd_sc_hd__mux2_1
XFILLER_101_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24801_ _10629_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25781_ _11180_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
X_34979_ clknet_leaf_472_CLK _03093_ VGND VGND VPWR VPWR registers\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_22993_ _09591_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27520_ _11822_ registers\[35\]\[44\] _12122_ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_444_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_444_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24732_ _10593_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21944_ registers\[52\]\[36\] registers\[53\]\[36\] registers\[54\]\[36\] registers\[55\]\[36\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__mux4_1
XFILLER_131_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27451_ _11753_ registers\[35\]\[11\] _12089_ VGND VGND VPWR VPWR _12091_ sky130_fd_sc_hd__mux2_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24663_ _09594_ registers\[55\]\[38\] _10547_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_24__f_CLK clknet_5_12_0_CLK VGND VGND VPWR VPWR clknet_6_24__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_21875_ _08326_ _08538_ _08539_ _08332_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__a22o_1
XFILLER_199_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26402_ _10852_ registers\[43\]\[58\] _11498_ VGND VGND VPWR VPWR _11507_ sky130_fd_sc_hd__mux2_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _09969_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20826_ registers\[4\]\[4\] registers\[5\]\[4\] registers\[6\]\[4\] registers\[7\]\[4\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__mux4_1
X_27382_ _12054_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__clkbuf_1
X_24594_ _09525_ registers\[55\]\[5\] _10514_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__mux2_1
XFILLER_70_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29121_ registers\[23\]\[22\] _12981_ _12977_ VGND VGND VPWR VPWR _12982_ sky130_fd_sc_hd__mux2_1
X_26333_ _10783_ registers\[43\]\[25\] _11465_ VGND VGND VPWR VPWR _11471_ sky130_fd_sc_hd__mux2_1
X_23545_ _09632_ registers\[19\]\[56\] _09925_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__mux2_1
X_20757_ registers\[0\]\[2\] registers\[1\]\[2\] registers\[2\]\[2\] registers\[3\]\[2\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__mux4_1
XFILLER_195_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29052_ _12934_ VGND VGND VPWR VPWR _12935_ sky130_fd_sc_hd__buf_4
XFILLER_195_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26264_ _11434_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
X_20688_ _07377_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__buf_6
X_23476_ _09563_ registers\[19\]\[23\] _09892_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__mux2_1
XFILLER_183_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28003_ _11763_ registers\[31\]\[16\] _12375_ VGND VGND VPWR VPWR _12382_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25215_ _10878_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__clkbuf_1
X_22427_ registers\[32\]\[50\] registers\[33\]\[50\] registers\[34\]\[50\] registers\[35\]\[50\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__mux4_1
XFILLER_137_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26195_ _11398_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25146_ net46 VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__buf_2
XFILLER_164_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22358_ registers\[36\]\[48\] registers\[37\]\[48\] registers\[38\]\[48\] registers\[39\]\[48\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__mux4_1
XFILLER_3_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21309_ _07983_ _07985_ _07988_ _07989_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__a22o_1
X_22289_ _08812_ _08940_ _08941_ _08815_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__a22o_1
XFILLER_3_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29954_ _13439_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__clkbuf_1
X_25077_ _10788_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28905_ _11855_ registers\[25\]\[60\] _12789_ VGND VGND VPWR VPWR _12856_ sky130_fd_sc_hd__mux2_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24028_ _10189_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29885_ registers\[18\]\[45\] _13029_ _13397_ VGND VGND VPWR VPWR _13403_ sky130_fd_sc_hd__mux2_1
XFILLER_133_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16850_ registers\[44\]\[22\] registers\[45\]\[22\] registers\[46\]\[22\] registers\[47\]\[22\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15342_ sky130_fd_sc_hd__mux4_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28836_ _11786_ registers\[25\]\[27\] _12812_ VGND VGND VPWR VPWR _12820_ sky130_fd_sc_hd__mux2_1
XFILLER_172_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28767_ _12783_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16781_ registers\[52\]\[20\] registers\[53\]\[20\] registers\[54\]\[20\] registers\[55\]\[20\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15275_ sky130_fd_sc_hd__mux4_1
X_25979_ _11284_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18520_ _05089_ _05277_ _05278_ _05100_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_435_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_435_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_218_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27718_ registers\[33\]\[9\] _10323_ _12222_ VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__mux2_1
XFILLER_19_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28698_ _12747_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__clkbuf_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18451_ _05077_ _05210_ _05211_ _05086_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a22o_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27649_ registers\[34\]\[40\] _10388_ _12195_ VGND VGND VPWR VPWR _12196_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_130 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_141 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ registers\[32\]\[38\] registers\[33\]\[38\] registers\[34\]\[38\] registers\[35\]\[38\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15878_ sky130_fd_sc_hd__mux4_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ registers\[16\]\[0\] registers\[17\]\[0\] registers\[18\]\[0\] registers\[19\]\[0\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__mux4_1
X_30660_ registers\[12\]\[28\] _12993_ _13802_ VGND VGND VPWR VPWR _13811_ sky130_fd_sc_hd__mux2_1
XANTENNA_163 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_196 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29319_ _13105_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__clkbuf_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _15677_ _15809_ _15810_ _15682_ VGND VGND VPWR VPWR _15811_ sky130_fd_sc_hd__a22o_1
XFILLER_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30591_ _13774_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__clkbuf_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32330_ clknet_leaf_152_CLK _00444_ VGND VGND VPWR VPWR registers\[19\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17264_ _15744_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19003_ _05080_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__clkbuf_4
X_16215_ registers\[48\]\[4\] registers\[49\]\[4\] registers\[50\]\[4\] registers\[51\]\[4\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14725_ sky130_fd_sc_hd__mux4_1
X_32261_ clknet_leaf_260_CLK _00375_ VGND VGND VPWR VPWR registers\[39\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_17195_ _14527_ VGND VGND VPWR VPWR _15677_ sky130_fd_sc_hd__buf_2
X_34000_ clknet_leaf_135_CLK _02114_ VGND VGND VPWR VPWR registers\[36\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31212_ _14101_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__clkbuf_1
X_16146_ _14581_ VGND VGND VPWR VPWR _14658_ sky130_fd_sc_hd__buf_6
XFILLER_128_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32192_ clknet_leaf_459_CLK _00306_ VGND VGND VPWR VPWR registers\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31143_ _14065_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__clkbuf_1
X_16077_ registers\[24\]\[0\] registers\[25\]\[0\] registers\[26\]\[0\] registers\[27\]\[0\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _14591_ sky130_fd_sc_hd__mux4_1
XFILLER_68_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19905_ registers\[12\]\[43\] registers\[13\]\[43\] registers\[14\]\[43\] registers\[15\]\[43\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__mux4_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35951_ clknet_leaf_378_CLK _04065_ VGND VGND VPWR VPWR registers\[6\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_31074_ registers\[0\]\[32\] _13002_ _14026_ VGND VGND VPWR VPWR _14029_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34902_ clknet_leaf_99_CLK _03016_ VGND VGND VPWR VPWR registers\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_30025_ _13476_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19836_ registers\[4\]\[41\] registers\[5\]\[41\] registers\[6\]\[41\] registers\[7\]\[41\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__mux4_1
XFILLER_233_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35882_ clknet_leaf_401_CLK _03996_ VGND VGND VPWR VPWR registers\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34833_ clknet_leaf_114_CLK _02947_ VGND VGND VPWR VPWR registers\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19767_ registers\[28\]\[39\] registers\[29\]\[39\] registers\[30\]\[39\] registers\[31\]\[39\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__mux4_1
Xinput3 DW[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_8
X_16979_ registers\[32\]\[26\] registers\[33\]\[26\] registers\[34\]\[26\] registers\[35\]\[26\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15467_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_426_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_426_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18718_ _05053_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__clkbuf_4
X_34764_ clknet_leaf_147_CLK _02878_ VGND VGND VPWR VPWR registers\[25\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_19698_ _06420_ _06423_ _06194_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__o21ba_1
X_31976_ clknet_leaf_6_CLK _00146_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
XFILLER_224_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33715_ clknet_leaf_346_CLK _01829_ VGND VGND VPWR VPWR registers\[41\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_782 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18649_ _05076_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__clkbuf_4
X_30927_ _13951_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__clkbuf_1
X_34695_ clknet_leaf_219_CLK _02809_ VGND VGND VPWR VPWR registers\[26\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30858_ _09815_ registers\[11\]\[58\] _13906_ VGND VGND VPWR VPWR _13915_ sky130_fd_sc_hd__mux2_1
XFILLER_197_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33646_ clknet_leaf_348_CLK _01760_ VGND VGND VPWR VPWR registers\[42\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_21660_ registers\[48\]\[28\] registers\[49\]\[28\] registers\[50\]\[28\] registers\[51\]\[28\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__mux4_1
XFILLER_80_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20611_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__buf_2
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21591_ registers\[52\]\[26\] registers\[53\]\[26\] registers\[54\]\[26\] registers\[55\]\[26\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__mux4_1
X_33577_ clknet_leaf_429_CLK _01691_ VGND VGND VPWR VPWR registers\[43\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_30789_ _09742_ registers\[11\]\[25\] _13873_ VGND VGND VPWR VPWR _13879_ sky130_fd_sc_hd__mux2_1
XFILLER_138_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20542_ _07239_ _07242_ _05162_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__o21ba_1
X_23330_ net54 VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__buf_4
X_35316_ clknet_leaf_416_CLK _03430_ VGND VGND VPWR VPWR registers\[16\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_824 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32528_ clknet_leaf_108_CLK _00642_ VGND VGND VPWR VPWR registers\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20473_ registers\[4\]\[60\] registers\[5\]\[60\] registers\[6\]\[60\] registers\[7\]\[60\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__mux4_1
X_35247_ clknet_leaf_394_CLK _03361_ VGND VGND VPWR VPWR registers\[17\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_23261_ net31 VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__clkbuf_4
X_32459_ clknet_leaf_158_CLK _00573_ VGND VGND VPWR VPWR registers\[29\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_25000_ _10736_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
X_22212_ registers\[28\]\[43\] registers\[29\]\[43\] registers\[30\]\[43\] registers\[31\]\[43\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__mux4_1
X_23192_ _09726_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35178_ clknet_leaf_406_CLK _03292_ VGND VGND VPWR VPWR registers\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22143_ registers\[20\]\[41\] registers\[21\]\[41\] registers\[22\]\[41\] registers\[23\]\[41\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__mux4_1
X_34129_ clknet_leaf_128_CLK _02243_ VGND VGND VPWR VPWR registers\[34\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26951_ _11816_ registers\[3\]\[41\] _11814_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__mux2_1
X_22074_ registers\[32\]\[40\] registers\[33\]\[40\] registers\[34\]\[40\] registers\[35\]\[40\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__mux4_1
XTAP_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21025_ registers\[48\]\[10\] registers\[49\]\[10\] registers\[50\]\[10\] registers\[51\]\[10\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__mux4_1
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25902_ _11244_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
X_29670_ registers\[1\]\[7\] _12949_ _13282_ VGND VGND VPWR VPWR _13290_ sky130_fd_sc_hd__mux2_1
X_26882_ _11769_ registers\[3\]\[19\] _11751_ VGND VGND VPWR VPWR _11770_ sky130_fd_sc_hd__mux2_1
XFILLER_102_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28621_ _11841_ registers\[27\]\[53\] _12703_ VGND VGND VPWR VPWR _12707_ sky130_fd_sc_hd__mux2_1
X_25833_ _10823_ registers\[47\]\[44\] _11203_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__mux2_1
XFILLER_68_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_417_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_417_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28552_ _11771_ registers\[27\]\[20\] _12670_ VGND VGND VPWR VPWR _12671_ sky130_fd_sc_hd__mux2_1
X_25764_ _10754_ registers\[47\]\[11\] _11170_ VGND VGND VPWR VPWR _11172_ sky130_fd_sc_hd__mux2_1
XFILLER_90_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22976_ net25 VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27503_ _11805_ registers\[35\]\[36\] _12111_ VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__mux2_1
XFILLER_56_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24715_ _09646_ registers\[55\]\[63\] _10513_ VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__mux2_1
XFILLER_15_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28483_ _12634_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21927_ _08423_ _08589_ _08590_ _08428_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__a22o_1
X_25695_ _11134_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27434_ _11736_ registers\[35\]\[3\] _12078_ VGND VGND VPWR VPWR _12082_ sky130_fd_sc_hd__mux2_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _10513_ VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21858_ _08418_ _08522_ _08523_ _08421_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__a22o_1
XFILLER_93_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20809_ registers\[44\]\[4\] registers\[45\]\[4\] registers\[46\]\[4\] registers\[47\]\[4\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__mux4_1
XFILLER_19_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27365_ _12045_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24577_ _09646_ registers\[56\]\[63\] _10439_ VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__mux2_1
XFILLER_24_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21789_ registers\[28\]\[31\] registers\[29\]\[31\] registers\[30\]\[31\] registers\[31\]\[31\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__mux4_1
X_29104_ net9 VGND VGND VPWR VPWR _12970_ sky130_fd_sc_hd__buf_2
XFILLER_204_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26316_ _10766_ registers\[43\]\[17\] _11454_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__mux2_1
XFILLER_184_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23528_ _09615_ registers\[19\]\[48\] _09914_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__mux2_1
XFILLER_243_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27296_ _12009_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29035_ _12924_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__clkbuf_1
X_26247_ _11425_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
X_23459_ _09546_ registers\[19\]\[15\] _09881_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__mux2_1
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16000_ registers\[44\]\[0\] registers\[45\]\[0\] registers\[46\]\[0\] registers\[47\]\[0\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14514_ sky130_fd_sc_hd__mux4_1
XFILLER_136_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26178_ _11389_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25129_ _10823_ registers\[52\]\[44\] _10815_ VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29937_ _13430_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__clkbuf_1
X_17951_ _04548_ _04723_ _04724_ _04552_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__a22o_1
XFILLER_174_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16902_ _15387_ _15392_ _15288_ VGND VGND VPWR VPWR _15393_ sky130_fd_sc_hd__o21ba_1
XFILLER_239_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17882_ registers\[52\]\[51\] registers\[53\]\[51\] registers\[54\]\[51\] registers\[55\]\[51\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__mux4_1
XFILLER_26_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29868_ registers\[18\]\[37\] _13012_ _13386_ VGND VGND VPWR VPWR _13394_ sky130_fd_sc_hd__mux2_1
XFILLER_215_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19621_ _06345_ _06348_ _06180_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__o21ba_1
X_28819_ _11769_ registers\[25\]\[19\] _12801_ VGND VGND VPWR VPWR _12811_ sky130_fd_sc_hd__mux2_1
X_16833_ registers\[24\]\[21\] registers\[25\]\[21\] registers\[26\]\[21\] registers\[27\]\[21\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15326_ sky130_fd_sc_hd__mux4_1
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29799_ registers\[18\]\[4\] _12943_ _13353_ VGND VGND VPWR VPWR _13358_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_408_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_408_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31830_ _14426_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19552_ registers\[12\]\[33\] registers\[13\]\[33\] registers\[14\]\[33\] registers\[15\]\[33\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__mux4_1
X_16764_ _15255_ _15258_ _14959_ VGND VGND VPWR VPWR _15259_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18503_ _05259_ _05262_ _05163_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__o21ba_1
XFILLER_74_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31761_ registers\[59\]\[38\] net32 _14381_ VGND VGND VPWR VPWR _14390_ sky130_fd_sc_hd__mux2_1
X_19483_ registers\[4\]\[31\] registers\[5\]\[31\] registers\[6\]\[31\] registers\[7\]\[31\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__mux4_1
X_16695_ registers\[40\]\[18\] registers\[41\]\[18\] registers\[42\]\[18\] registers\[43\]\[18\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15191_ sky130_fd_sc_hd__mux4_1
XFILLER_34_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30712_ _13838_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__clkbuf_1
X_33500_ clknet_leaf_30_CLK _01614_ VGND VGND VPWR VPWR registers\[44\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18434_ _05174_ _05181_ _05188_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__or4_4
XFILLER_146_1227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31692_ registers\[59\]\[5\] net56 _14348_ VGND VGND VPWR VPWR _14354_ sky130_fd_sc_hd__mux2_1
XFILLER_22_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34480_ clknet_leaf_377_CLK _02594_ VGND VGND VPWR VPWR registers\[2\]\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_871 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33431_ clknet_leaf_123_CLK _01545_ VGND VGND VPWR VPWR registers\[45\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_18365_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30643_ _13779_ VGND VGND VPWR VPWR _13802_ sky130_fd_sc_hd__buf_4
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17316_ registers\[0\]\[35\] registers\[1\]\[35\] registers\[2\]\[35\] registers\[3\]\[35\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15795_ sky130_fd_sc_hd__mux4_1
X_33362_ clknet_leaf_123_CLK _01476_ VGND VGND VPWR VPWR registers\[46\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_36150_ clknet_leaf_335_CLK _04264_ VGND VGND VPWR VPWR registers\[49\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_30574_ _09800_ registers\[13\]\[51\] _13764_ VGND VGND VPWR VPWR _13766_ sky130_fd_sc_hd__mux2_1
X_18296_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__buf_12
X_35101_ clknet_leaf_478_CLK _03215_ VGND VGND VPWR VPWR registers\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_32313_ clknet_leaf_309_CLK _00427_ VGND VGND VPWR VPWR registers\[19\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17247_ registers\[8\]\[33\] registers\[9\]\[33\] registers\[10\]\[33\] registers\[11\]\[33\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15728_ sky130_fd_sc_hd__mux4_1
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33293_ clknet_leaf_169_CLK _01407_ VGND VGND VPWR VPWR registers\[48\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_36081_ clknet_leaf_366_CLK _04195_ VGND VGND VPWR VPWR registers\[59\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_35032_ clknet_leaf_487_CLK _03146_ VGND VGND VPWR VPWR registers\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_32244_ clknet_leaf_350_CLK _00358_ VGND VGND VPWR VPWR registers\[39\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_17178_ _15657_ _15660_ _15620_ _15621_ VGND VGND VPWR VPWR _15661_ sky130_fd_sc_hd__o211a_1
XFILLER_115_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ _14588_ _14640_ _14641_ _14598_ VGND VGND VPWR VPWR _14642_ sky130_fd_sc_hd__a22o_1
X_32175_ clknet_leaf_12_CLK _00289_ VGND VGND VPWR VPWR registers\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31126_ registers\[0\]\[57\] _13054_ _14048_ VGND VGND VPWR VPWR _14056_ sky130_fd_sc_hd__mux2_1
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35934_ clknet_leaf_481_CLK _04048_ VGND VGND VPWR VPWR registers\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31057_ registers\[0\]\[24\] _12985_ _14015_ VGND VGND VPWR VPWR _14020_ sky130_fd_sc_hd__mux2_1
XFILLER_243_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30008_ _13467_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19819_ registers\[32\]\[41\] registers\[33\]\[41\] registers\[34\]\[41\] registers\[35\]\[41\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__mux4_1
X_35865_ clknet_leaf_475_CLK _03979_ VGND VGND VPWR VPWR registers\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34816_ clknet_leaf_225_CLK _02930_ VGND VGND VPWR VPWR registers\[24\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_22830_ registers\[0\]\[62\] registers\[1\]\[62\] registers\[2\]\[62\] registers\[3\]\[62\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__mux4_1
XFILLER_238_891 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35796_ clknet_leaf_81_CLK _03910_ VGND VGND VPWR VPWR registers\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22761_ _09396_ _09399_ _07309_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__o21ba_1
X_34747_ clknet_leaf_187_CLK _02861_ VGND VGND VPWR VPWR registers\[25\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_213_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31959_ clknet_leaf_0_CLK _00191_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_1
X_24500_ _09569_ registers\[56\]\[26\] _10462_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__mux2_1
XFILLER_240_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21712_ registers\[16\]\[29\] registers\[17\]\[29\] registers\[18\]\[29\] registers\[19\]\[29\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__mux4_1
X_25480_ registers\[4\]\[7\] _10319_ _11012_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22692_ _09330_ _09333_ _09116_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34678_ clknet_leaf_312_CLK _02792_ VGND VGND VPWR VPWR registers\[26\]\[40\] sky130_fd_sc_hd__dfxtp_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24431_ net57 VGND VGND VPWR VPWR _10430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_240_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21643_ registers\[20\]\[27\] registers\[21\]\[27\] registers\[22\]\[27\] registers\[23\]\[27\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__mux4_1
X_33629_ clknet_leaf_28_CLK _01743_ VGND VGND VPWR VPWR registers\[42\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27150_ _11857_ registers\[38\]\[61\] _11864_ VGND VGND VPWR VPWR _11932_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24362_ _10383_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_30 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21574_ _08080_ _08246_ _08247_ _08085_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__a22o_1
XFILLER_205_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_41 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26101_ _10821_ registers\[45\]\[43\] _11345_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__mux2_1
X_23313_ net49 VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__buf_4
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_63 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20525_ registers\[60\]\[62\] registers\[61\]\[62\] registers\[62\]\[62\] registers\[63\]\[62\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__mux4_1
X_27081_ _11788_ registers\[38\]\[28\] _11887_ VGND VGND VPWR VPWR _11896_ sky130_fd_sc_hd__mux2_1
XANTENNA_74 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24293_ registers\[57\]\[15\] _10336_ _10326_ VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__mux2_1
XANTENNA_85 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26032_ _10751_ registers\[45\]\[10\] _11312_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__mux2_1
XFILLER_107_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20456_ registers\[32\]\[60\] registers\[33\]\[60\] registers\[34\]\[60\] registers\[35\]\[60\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__mux4_1
XFILLER_153_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23244_ net26 VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20387_ registers\[16\]\[57\] registers\[17\]\[57\] registers\[18\]\[57\] registers\[19\]\[57\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__mux4_2
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23175_ net15 VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22126_ registers\[48\]\[41\] registers\[49\]\[41\] registers\[50\]\[41\] registers\[51\]\[41\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__mux4_1
XANTENNA_1309 _00150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27983_ _12371_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__clkbuf_1
XTAP_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput170 net170 VGND VGND VPWR VPWR D2[24] sky130_fd_sc_hd__buf_2
XTAP_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput181 net181 VGND VGND VPWR VPWR D2[34] sky130_fd_sc_hd__buf_2
XTAP_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput192 net192 VGND VGND VPWR VPWR D2[44] sky130_fd_sc_hd__buf_2
XTAP_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29722_ _13317_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__clkbuf_1
X_26934_ net30 VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22057_ registers\[8\]\[39\] registers\[9\]\[39\] registers\[10\]\[39\] registers\[11\]\[39\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__mux4_1
XFILLER_212_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ registers\[28\]\[9\] registers\[29\]\[9\] registers\[30\]\[9\] registers\[31\]\[9\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__mux4_1
XFILLER_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29653_ _13280_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__clkbuf_1
XTAP_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26865_ _11758_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_1
XTAP_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28604_ _11824_ registers\[27\]\[45\] _12692_ VGND VGND VPWR VPWR _12698_ sky130_fd_sc_hd__mux2_1
X_25816_ _10806_ registers\[47\]\[36\] _11192_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__mux2_1
X_29584_ registers\[20\]\[30\] _12997_ _13244_ VGND VGND VPWR VPWR _13245_ sky130_fd_sc_hd__mux2_1
X_26796_ _11715_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28535_ _11755_ registers\[27\]\[12\] _12659_ VGND VGND VPWR VPWR _12662_ sky130_fd_sc_hd__mux2_1
X_25747_ _10737_ registers\[47\]\[3\] _11159_ VGND VGND VPWR VPWR _11163_ sky130_fd_sc_hd__mux2_1
XFILLER_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22959_ _09568_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28466_ _12625_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ registers\[24\]\[11\] registers\[25\]\[11\] registers\[26\]\[11\] registers\[27\]\[11\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14983_ sky130_fd_sc_hd__mux4_1
XFILLER_189_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25678_ _11125_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27417_ _12072_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24629_ _10538_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28397_ _12589_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__clkbuf_1
X_18150_ registers\[20\]\[59\] registers\[21\]\[59\] registers\[22\]\[59\] registers\[23\]\[59\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__mux4_1
XFILLER_175_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27348_ _12036_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17101_ registers\[52\]\[29\] registers\[53\]\[29\] registers\[54\]\[29\] registers\[55\]\[29\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15586_ sky130_fd_sc_hd__mux4_1
XFILLER_15_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18081_ _14491_ _04849_ _04850_ _14501_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a22o_1
XFILLER_89_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27279_ _11851_ registers\[37\]\[58\] _11991_ VGND VGND VPWR VPWR _12000_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29018_ _12915_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__clkbuf_1
X_17032_ registers\[8\]\[27\] registers\[9\]\[27\] registers\[10\]\[27\] registers\[11\]\[27\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15519_ sky130_fd_sc_hd__mux4_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30290_ registers\[15\]\[45\] _13029_ _13610_ VGND VGND VPWR VPWR _13616_ sky130_fd_sc_hd__mux2_1
XFILLER_194_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ registers\[4\]\[17\] registers\[5\]\[17\] registers\[6\]\[17\] registers\[7\]\[17\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__mux4_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ registers\[20\]\[52\] registers\[21\]\[52\] registers\[22\]\[52\] registers\[23\]\[52\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__mux4_1
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33980_ clknet_leaf_276_CLK _02094_ VGND VGND VPWR VPWR registers\[37\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32931_ clknet_leaf_443_CLK _01045_ VGND VGND VPWR VPWR registers\[53\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17865_ _14581_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19604_ _06233_ _06330_ _06331_ _06236_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__a22o_1
X_35650_ clknet_leaf_242_CLK _03764_ VGND VGND VPWR VPWR registers\[11\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_16816_ registers\[36\]\[21\] registers\[37\]\[21\] registers\[38\]\[21\] registers\[39\]\[21\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15309_ sky130_fd_sc_hd__mux4_1
X_32862_ clknet_leaf_46_CLK _00976_ VGND VGND VPWR VPWR registers\[54\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_17796_ _14504_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__buf_4
XFILLER_213_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34601_ clknet_leaf_453_CLK _02715_ VGND VGND VPWR VPWR registers\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31813_ registers\[59\]\[63\] net60 _14347_ VGND VGND VPWR VPWR _14417_ sky130_fd_sc_hd__mux2_1
X_19535_ _06226_ _06263_ _06264_ _06231_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a22o_1
X_35581_ clknet_leaf_297_CLK _03695_ VGND VGND VPWR VPWR registers\[12\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_16747_ registers\[60\]\[19\] registers\[61\]\[19\] registers\[62\]\[19\] registers\[63\]\[19\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15242_ sky130_fd_sc_hd__mux4_1
X_32793_ clknet_leaf_66_CLK _00907_ VGND VGND VPWR VPWR registers\[55\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34532_ clknet_leaf_464_CLK _02646_ VGND VGND VPWR VPWR registers\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31744_ _14347_ VGND VGND VPWR VPWR _14381_ sky130_fd_sc_hd__buf_4
X_19466_ registers\[32\]\[31\] registers\[33\]\[31\] registers\[34\]\[31\] registers\[35\]\[31\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__mux4_1
X_16678_ _15171_ _15174_ _14934_ _14935_ VGND VGND VPWR VPWR _15175_ sky130_fd_sc_hd__o211a_1
XFILLER_222_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18417_ registers\[52\]\[1\] registers\[53\]\[1\] registers\[54\]\[1\] registers\[55\]\[1\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__mux4_1
XFILLER_50_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34463_ clknet_leaf_487_CLK _02577_ VGND VGND VPWR VPWR registers\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_31675_ _14344_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19397_ registers\[56\]\[29\] registers\[57\]\[29\] registers\[58\]\[29\] registers\[59\]\[29\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux4_1
X_36202_ clknet_leaf_92_CLK _00084_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dfxtp_1
X_33414_ clknet_leaf_254_CLK _01528_ VGND VGND VPWR VPWR registers\[46\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_18348_ _05078_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__buf_12
X_30626_ _13793_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__clkbuf_1
X_34394_ clknet_leaf_4_CLK _02508_ VGND VGND VPWR VPWR registers\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36133_ clknet_leaf_440_CLK _04247_ VGND VGND VPWR VPWR registers\[49\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_33345_ clknet_leaf_258_CLK _01459_ VGND VGND VPWR VPWR registers\[47\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_18279_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__buf_12
X_30557_ _09782_ registers\[13\]\[43\] _13753_ VGND VGND VPWR VPWR _13757_ sky130_fd_sc_hd__mux2_1
XFILLER_124_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20310_ _06919_ _07016_ _07017_ _06922_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__a22o_1
XFILLER_174_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21290_ registers\[20\]\[17\] registers\[21\]\[17\] registers\[22\]\[17\] registers\[23\]\[17\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__mux4_1
Xinput50 DW[54] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_8
X_36064_ clknet_leaf_43_CLK _04178_ VGND VGND VPWR VPWR registers\[59\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33276_ clknet_leaf_276_CLK _01390_ VGND VGND VPWR VPWR registers\[48\]\[46\] sky130_fd_sc_hd__dfxtp_1
Xinput61 DW[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_6
X_30488_ _09678_ registers\[13\]\[10\] _13720_ VGND VGND VPWR VPWR _13721_ sky130_fd_sc_hd__mux2_1
Xinput72 R2[1] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput83 RW[0] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_4
X_20241_ _06912_ _06949_ _06950_ _06917_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__a22o_1
X_35015_ clknet_leaf_206_CLK _03129_ VGND VGND VPWR VPWR registers\[21\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_32227_ clknet_leaf_216_CLK _00341_ VGND VGND VPWR VPWR registers\[9\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20172_ registers\[32\]\[51\] registers\[33\]\[51\] registers\[34\]\[51\] registers\[35\]\[51\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux4_1
X_32158_ clknet_leaf_23_CLK _00272_ VGND VGND VPWR VPWR registers\[39\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1055 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31109_ registers\[0\]\[49\] _13037_ _14037_ VGND VGND VPWR VPWR _14047_ sky130_fd_sc_hd__mux2_1
X_24980_ _10723_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32089_ clknet_leaf_489_CLK _00002_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35917_ clknet_leaf_144_CLK _04031_ VGND VGND VPWR VPWR registers\[7\]\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ _09607_ registers\[60\]\[44\] _10133_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__mux2_1
XFILLER_229_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26650_ _10829_ registers\[41\]\[47\] _11630_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__mux2_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35848_ clknet_leaf_154_CLK _03962_ VGND VGND VPWR VPWR registers\[8\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_23862_ _09538_ registers\[60\]\[11\] _10100_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__mux2_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25601_ _11083_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22813_ _09429_ _09436_ _09443_ _09450_ VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__or4_4
XANTENNA_707 _07289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26581_ _10760_ registers\[41\]\[14\] _11597_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__mux2_1
X_35779_ clknet_leaf_241_CLK _03893_ VGND VGND VPWR VPWR registers\[0\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23793_ _09605_ registers\[29\]\[43\] _10061_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__mux2_1
XANTENNA_718 _07315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_729 _07352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28320_ _12548_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__clkbuf_1
X_25532_ _11047_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_1
X_22744_ _07296_ _09382_ _09383_ _07302_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__a22o_1
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28251_ _12512_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25463_ _11009_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__buf_6
XFILLER_198_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22675_ registers\[60\]\[57\] registers\[61\]\[57\] registers\[62\]\[57\] registers\[63\]\[57\]
+ _09227_ _09021_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__mux4_1
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27202_ _11774_ registers\[37\]\[21\] _11958_ VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__mux2_1
X_24414_ registers\[57\]\[54\] _10418_ _10410_ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28182_ _11807_ registers\[30\]\[37\] _12468_ VGND VGND VPWR VPWR _12476_ sky130_fd_sc_hd__mux2_1
X_21626_ registers\[48\]\[27\] registers\[49\]\[27\] registers\[50\]\[27\] registers\[51\]\[27\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__mux4_1
XFILLER_90_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25394_ _10798_ registers\[50\]\[32\] _10970_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__mux2_1
XFILLER_138_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27133_ _11923_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24345_ net26 VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__buf_4
XFILLER_138_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21557_ registers\[52\]\[25\] registers\[53\]\[25\] registers\[54\]\[25\] registers\[55\]\[25\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__mux4_1
XFILLER_240_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20508_ _05107_ _07208_ _07209_ _05117_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__a22o_1
X_27064_ _11864_ VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__buf_4
XFILLER_154_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24276_ net2 VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__buf_4
XFILLER_107_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21488_ registers\[48\]\[23\] registers\[49\]\[23\] registers\[50\]\[23\] registers\[51\]\[23\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__mux4_1
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26015_ _10735_ registers\[45\]\[2\] _11301_ VGND VGND VPWR VPWR _11304_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23227_ _09746_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
XTAP_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20439_ registers\[8\]\[59\] registers\[9\]\[59\] registers\[10\]\[59\] registers\[11\]\[59\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__mux4_1
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23158_ _09706_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__buf_6
XTAP_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1106 _14553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1117 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22109_ _07315_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__buf_4
XFILLER_121_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1128 _14600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15980_ _14493_ VGND VGND VPWR VPWR _14494_ sky130_fd_sc_hd__buf_6
X_23089_ _09659_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__clkbuf_1
XTAP_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1139 _14613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27966_ registers\[32\]\[63\] _10436_ _12292_ VGND VGND VPWR VPWR _12362_ sky130_fd_sc_hd__mux2_1
XTAP_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29705_ _13308_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26917_ _11792_ registers\[3\]\[30\] _11793_ VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__mux2_1
XTAP_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27897_ _12292_ VGND VGND VPWR VPWR _12326_ sky130_fd_sc_hd__buf_4
XTAP_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29636_ registers\[20\]\[55\] _13050_ _13266_ VGND VGND VPWR VPWR _13272_ sky130_fd_sc_hd__mux2_1
XTAP_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _04407_ _04416_ _04423_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__or4_2
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26848_ _11746_ registers\[3\]\[8\] _11730_ VGND VGND VPWR VPWR _11747_ sky130_fd_sc_hd__mux2_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ registers\[48\]\[15\] registers\[49\]\[15\] registers\[50\]\[15\] registers\[51\]\[15\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15100_ sky130_fd_sc_hd__mux4_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ registers\[20\]\[42\] registers\[21\]\[42\] registers\[22\]\[42\] registers\[23\]\[42\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__mux4_1
XFILLER_95_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26779_ _11706_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__clkbuf_1
X_29567_ registers\[20\]\[22\] _12981_ _13233_ VGND VGND VPWR VPWR _13236_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16532_ _14998_ _15031_ _15032_ _15001_ VGND VGND VPWR VPWR _15033_ sky130_fd_sc_hd__a22o_1
X_19320_ _05120_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__buf_6
XFILLER_186_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28518_ _11738_ registers\[27\]\[4\] _12648_ VGND VGND VPWR VPWR _12653_ sky130_fd_sc_hd__mux2_1
XFILLER_204_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29498_ _13199_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16463_ registers\[36\]\[11\] registers\[37\]\[11\] registers\[38\]\[11\] registers\[39\]\[11\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _14966_ sky130_fd_sc_hd__mux4_1
XFILLER_108_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19251_ _05890_ _05987_ _05988_ _05893_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__a22o_1
XFILLER_182_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28449_ _12616_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18202_ registers\[12\]\[61\] registers\[13\]\[61\] registers\[14\]\[61\] registers\[15\]\[61\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__mux4_1
XFILLER_204_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31460_ _09730_ registers\[6\]\[23\] _14228_ VGND VGND VPWR VPWR _14232_ sky130_fd_sc_hd__mux2_1
X_19182_ _05883_ _05920_ _05921_ _05888_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__a22o_1
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16394_ registers\[60\]\[9\] registers\[61\]\[9\] registers\[62\]\[9\] registers\[63\]\[9\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _14899_ sky130_fd_sc_hd__mux4_1
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ registers\[48\]\[59\] registers\[49\]\[59\] registers\[50\]\[59\] registers\[51\]\[59\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__mux4_1
X_30411_ _09771_ registers\[14\]\[38\] _13671_ VGND VGND VPWR VPWR _13680_ sky130_fd_sc_hd__mux2_1
XFILLER_8_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31391_ _14195_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_805 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18064_ _04834_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_2
X_30342_ _09668_ registers\[14\]\[5\] _13638_ VGND VGND VPWR VPWR _13644_ sky130_fd_sc_hd__mux2_1
X_33130_ clknet_leaf_420_CLK _01244_ VGND VGND VPWR VPWR registers\[50\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17015_ _15502_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33061_ clknet_leaf_440_CLK _01175_ VGND VGND VPWR VPWR registers\[51\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_30273_ registers\[15\]\[37\] _13012_ _13599_ VGND VGND VPWR VPWR _13607_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32012_ clknet_leaf_29_CLK _00186_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_1
XFILLER_171_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18966_ registers\[44\]\[17\] registers\[45\]\[17\] registers\[46\]\[17\] registers\[47\]\[17\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__mux4_1
XFILLER_239_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1640 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1651 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1662 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17917_ registers\[60\]\[52\] registers\[61\]\[52\] registers\[62\]\[52\] registers\[63\]\[52\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux4_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1673 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33963_ clknet_leaf_424_CLK _02077_ VGND VGND VPWR VPWR registers\[37\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_18897_ registers\[36\]\[15\] registers\[37\]\[15\] registers\[38\]\[15\] registers\[39\]\[15\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__mux4_1
XFILLER_239_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1684 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1695 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35702_ clknet_leaf_331_CLK _03816_ VGND VGND VPWR VPWR registers\[10\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_32914_ clknet_leaf_181_CLK _01028_ VGND VGND VPWR VPWR registers\[53\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17848_ registers\[0\]\[50\] registers\[1\]\[50\] registers\[2\]\[50\] registers\[3\]\[50\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__mux4_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33894_ clknet_leaf_433_CLK _02008_ VGND VGND VPWR VPWR registers\[38\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35633_ clknet_leaf_381_CLK _03747_ VGND VGND VPWR VPWR registers\[11\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_32845_ clknet_leaf_141_CLK _00959_ VGND VGND VPWR VPWR registers\[55\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_17779_ registers\[12\]\[48\] registers\[13\]\[48\] registers\[14\]\[48\] registers\[15\]\[48\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux4_1
XFILLER_240_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19518_ registers\[12\]\[32\] registers\[13\]\[32\] registers\[14\]\[32\] registers\[15\]\[32\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux4_1
XFILLER_241_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35564_ clknet_leaf_392_CLK _03678_ VGND VGND VPWR VPWR registers\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20790_ _07343_ _07484_ _07485_ _07353_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a22o_1
X_32776_ clknet_leaf_192_CLK _00890_ VGND VGND VPWR VPWR registers\[56\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34515_ clknet_leaf_103_CLK _02629_ VGND VGND VPWR VPWR registers\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19449_ _05136_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__clkbuf_4
X_31727_ _14372_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__clkbuf_1
X_35495_ clknet_leaf_460_CLK _03609_ VGND VGND VPWR VPWR registers\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22460_ _07295_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__clkbuf_4
X_34446_ clknet_leaf_109_CLK _02560_ VGND VGND VPWR VPWR registers\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31658_ registers\[63\]\[53\] net49 _14332_ VGND VGND VPWR VPWR _14336_ sky130_fd_sc_hd__mux2_1
XFILLER_163_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21411_ _08089_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30609_ _13784_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__clkbuf_1
X_34377_ clknet_leaf_214_CLK _02491_ VGND VGND VPWR VPWR registers\[31\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_22391_ _09038_ _09041_ _08773_ VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__o21ba_1
XFILLER_241_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31589_ registers\[63\]\[20\] net13 _14299_ VGND VGND VPWR VPWR _14300_ sky130_fd_sc_hd__mux2_1
XFILLER_108_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36116_ clknet_leaf_70_CLK _04230_ VGND VGND VPWR VPWR registers\[49\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_24130_ _10243_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33328_ clknet_leaf_362_CLK _01442_ VGND VGND VPWR VPWR registers\[47\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_21342_ _07783_ _08020_ _08021_ _07786_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__a22o_1
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36047_ clknet_leaf_173_CLK _04161_ VGND VGND VPWR VPWR registers\[59\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_24061_ _09601_ registers\[5\]\[41\] _10205_ VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__mux2_1
X_21273_ registers\[48\]\[17\] registers\[49\]\[17\] registers\[50\]\[17\] registers\[51\]\[17\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__mux4_1
X_33259_ clknet_leaf_425_CLK _01373_ VGND VGND VPWR VPWR registers\[48\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23012_ _09604_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20224_ registers\[12\]\[52\] registers\[13\]\[52\] registers\[14\]\[52\] registers\[15\]\[52\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__mux4_1
XFILLER_46_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27820_ _12285_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__clkbuf_1
X_20155_ _05039_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24963_ _09622_ registers\[53\]\[51\] _10713_ VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__mux2_1
X_20086_ registers\[16\]\[48\] registers\[17\]\[48\] registers\[18\]\[48\] registers\[19\]\[48\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__mux4_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27751_ _12249_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__clkbuf_1
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26702_ registers\[40\]\[7\] _10319_ _11658_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23914_ _09590_ registers\[60\]\[36\] _10122_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__mux2_1
X_27682_ registers\[34\]\[56\] _10422_ _12206_ VGND VGND VPWR VPWR _12213_ sky130_fd_sc_hd__mux2_1
XFILLER_217_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24894_ _10678_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29421_ _09693_ registers\[21\]\[17\] _13151_ VGND VGND VPWR VPWR _13159_ sky130_fd_sc_hd__mux2_1
XFILLER_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26633_ _10812_ registers\[41\]\[39\] _11619_ VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__mux2_1
X_23845_ _09521_ registers\[60\]\[3\] _10089_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__mux2_1
XFILLER_150_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_504 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_515 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_526 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_537 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26564_ _10743_ registers\[41\]\[6\] _11586_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__mux2_1
X_29352_ _13122_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__clkbuf_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_548 _04352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23776_ _09588_ registers\[29\]\[35\] _10050_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__mux2_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20988_ registers\[36\]\[9\] registers\[37\]\[9\] registers\[38\]\[9\] registers\[39\]\[9\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__mux4_1
XANTENNA_559 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25515_ _11038_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__clkbuf_1
X_28303_ registers\[2\]\[30\] _10367_ _12539_ VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__mux2_1
X_22727_ _09148_ _09365_ _09366_ _09153_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__a22o_1
X_29283_ _13086_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_886 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26495_ _10810_ registers\[42\]\[38\] _11547_ VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28234_ _11859_ registers\[30\]\[62\] _12434_ VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__mux2_1
X_25446_ _10850_ registers\[50\]\[57\] _10992_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__mux2_1
X_22658_ _09104_ _09299_ _09300_ _09107_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__a22o_1
XFILLER_139_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28165_ _11790_ registers\[30\]\[29\] _12457_ VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__mux2_1
X_21609_ _08075_ _08278_ _08281_ _08078_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__a22o_1
X_25377_ _10781_ registers\[50\]\[24\] _10959_ VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__mux2_1
X_22589_ _08953_ _09232_ _09233_ _08956_ VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__a22o_1
XFILLER_220_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27116_ _11914_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24328_ _10360_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
X_28096_ _12430_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27047_ _11878_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__clkbuf_1
X_24259_ registers\[57\]\[4\] _10313_ _10305_ VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__mux2_1
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18820_ _05152_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__buf_4
XTAP_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1056 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28998_ net282 VGND VGND VPWR VPWR _12905_ sky130_fd_sc_hd__buf_4
XTAP_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18751_ _05156_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__buf_4
X_27949_ _12353_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__clkbuf_1
XTAP_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ registers\[0\]\[46\] registers\[1\]\[46\] registers\[2\]\[46\] registers\[3\]\[46\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__mux4_1
XFILLER_208_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18682_ registers\[40\]\[9\] registers\[41\]\[9\] registers\[42\]\[9\] registers\[43\]\[9\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__mux4_1
XTAP_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30960_ registers\[10\]\[42\] _13023_ _13966_ VGND VGND VPWR VPWR _13969_ sky130_fd_sc_hd__mux2_1
XTAP_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29619_ registers\[20\]\[47\] _13033_ _13255_ VGND VGND VPWR VPWR _13263_ sky130_fd_sc_hd__mux2_1
X_17633_ _04411_ _04415_ _15963_ _15964_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__o211a_1
XFILLER_64_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30891_ _13932_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32630_ clknet_leaf_329_CLK _00744_ VGND VGND VPWR VPWR registers\[58\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_17564_ registers\[60\]\[42\] registers\[61\]\[42\] registers\[62\]\[42\] registers\[63\]\[42\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__mux4_1
XFILLER_216_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19303_ _06036_ _06037_ _06038_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__a22o_1
XFILLER_32_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16515_ _15013_ _15016_ _14945_ VGND VGND VPWR VPWR _15017_ sky130_fd_sc_hd__o21ba_1
XFILLER_225_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32561_ clknet_leaf_372_CLK _00675_ VGND VGND VPWR VPWR registers\[5\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ registers\[0\]\[40\] registers\[1\]\[40\] registers\[2\]\[40\] registers\[3\]\[40\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _15969_ sky130_fd_sc_hd__mux4_1
X_34300_ clknet_leaf_277_CLK _02414_ VGND VGND VPWR VPWR registers\[32\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_31512_ _09793_ registers\[6\]\[48\] _14250_ VGND VGND VPWR VPWR _14259_ sky130_fd_sc_hd__mux2_1
X_19234_ _05969_ _05972_ _05837_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35280_ clknet_leaf_112_CLK _03394_ VGND VGND VPWR VPWR registers\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16446_ _14597_ VGND VGND VPWR VPWR _14950_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32492_ clknet_leaf_370_CLK _00606_ VGND VGND VPWR VPWR registers\[60\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34231_ clknet_leaf_342_CLK _02345_ VGND VGND VPWR VPWR registers\[33\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_16377_ registers\[20\]\[8\] registers\[21\]\[8\] registers\[22\]\[8\] registers\[23\]\[8\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14883_ sky130_fd_sc_hd__mux4_1
X_19165_ registers\[12\]\[22\] registers\[13\]\[22\] registers\[14\]\[22\] registers\[15\]\[22\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__mux4_1
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31443_ _09689_ registers\[6\]\[15\] _14217_ VGND VGND VPWR VPWR _14223_ sky130_fd_sc_hd__mux2_1
XFILLER_219_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18116_ registers\[24\]\[58\] registers\[25\]\[58\] registers\[26\]\[58\] registers\[27\]\[58\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__mux4_1
X_31374_ _14186_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34162_ clknet_leaf_359_CLK _02276_ VGND VGND VPWR VPWR registers\[34\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19096_ _05136_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__clkbuf_4
XFILLER_195_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30325_ registers\[15\]\[62\] _13064_ _13565_ VGND VGND VPWR VPWR _13634_ sky130_fd_sc_hd__mux2_1
X_33113_ clknet_leaf_84_CLK _01227_ VGND VGND VPWR VPWR registers\[50\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18047_ _04548_ _04816_ _04817_ _04552_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a22o_1
X_34093_ clknet_leaf_321_CLK _02207_ VGND VGND VPWR VPWR registers\[35\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33044_ clknet_leaf_70_CLK _01158_ VGND VGND VPWR VPWR registers\[51\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30256_ registers\[15\]\[29\] _12995_ _13588_ VGND VGND VPWR VPWR _13598_ sky130_fd_sc_hd__mux2_1
XFILLER_236_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30187_ _13561_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19998_ _06441_ _06711_ _06714_ _06445_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__a22o_1
XFILLER_45_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18949_ _05130_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__clkbuf_4
X_34995_ clknet_leaf_384_CLK _03109_ VGND VGND VPWR VPWR registers\[21\]\[37\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1470 _05328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1481 _06051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1492 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21960_ _07317_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__buf_4
X_33946_ clknet_leaf_22_CLK _02060_ VGND VGND VPWR VPWR registers\[37\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20911_ registers\[32\]\[7\] registers\[33\]\[7\] registers\[34\]\[7\] registers\[35\]\[7\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__mux4_1
XFILLER_243_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33877_ clknet_leaf_117_CLK _01991_ VGND VGND VPWR VPWR registers\[38\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_21891_ registers\[16\]\[34\] registers\[17\]\[34\] registers\[18\]\[34\] registers\[19\]\[34\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__mux4_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35616_ clknet_leaf_485_CLK _03730_ VGND VGND VPWR VPWR registers\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_23630_ registers\[61\]\[31\] _09756_ _09976_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__mux2_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20842_ _07433_ _07534_ _07535_ _07438_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__a22o_1
X_32828_ clknet_leaf_292_CLK _00942_ VGND VGND VPWR VPWR registers\[55\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_23561_ net83 _09512_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__nand2_8
X_35547_ clknet_leaf_477_CLK _03661_ VGND VGND VPWR VPWR registers\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_20773_ _07469_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32759_ clknet_leaf_328_CLK _00873_ VGND VGND VPWR VPWR registers\[56\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25300_ _10840_ registers\[51\]\[52\] _10920_ VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__mux2_1
XFILLER_211_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22512_ _09155_ _09156_ _09157_ _09158_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__a22o_1
X_26280_ _11442_ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__buf_4
XFILLER_222_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35478_ clknet_leaf_82_CLK _03592_ VGND VGND VPWR VPWR registers\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_23492_ _09904_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_867 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25231_ _10886_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22443_ _07340_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__clkbuf_4
X_34429_ clknet_leaf_183_CLK _02543_ VGND VGND VPWR VPWR registers\[30\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25162_ net51 VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__buf_2
XFILLER_176_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22374_ _09020_ _09022_ _09023_ _09024_ VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__a22o_1
XFILLER_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24113_ _09517_ registers\[58\]\[1\] _10233_ VGND VGND VPWR VPWR _10235_ sky130_fd_sc_hd__mux2_1
X_21325_ _08000_ _08005_ _07730_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__o21ba_1
X_25093_ _10799_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_1
X_29970_ registers\[17\]\[21\] _12979_ _13446_ VGND VGND VPWR VPWR _13448_ sky130_fd_sc_hd__mux2_1
XFILLER_190_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28921_ registers\[24\]\[3\] _10311_ _12861_ VGND VGND VPWR VPWR _12865_ sky130_fd_sc_hd__mux2_1
X_24044_ _09584_ registers\[5\]\[33\] _10194_ VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__mux2_1
X_21256_ _07732_ _07935_ _07938_ _07735_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__a22o_1
XFILLER_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_47__f_CLK clknet_5_23_0_CLK VGND VGND VPWR VPWR clknet_6_47__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20207_ _06912_ _06915_ _06916_ _06917_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__a22o_1
X_28852_ _12828_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__clkbuf_1
X_21187_ registers\[28\]\[14\] registers\[29\]\[14\] registers\[30\]\[14\] registers\[31\]\[14\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__mux4_1
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27803_ _12276_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__clkbuf_1
X_20138_ _06776_ _06849_ _06850_ _06782_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__a22o_1
X_25995_ _10850_ registers\[46\]\[57\] _11285_ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__mux2_1
X_28783_ _12792_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__clkbuf_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _05058_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__buf_4
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24946_ _09605_ registers\[53\]\[43\] _10702_ VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__mux2_1
X_27734_ _12240_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_1
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27665_ registers\[34\]\[48\] _10405_ _12195_ VGND VGND VPWR VPWR _12204_ sky130_fd_sc_hd__mux2_1
X_24877_ _09535_ registers\[53\]\[10\] _10669_ VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__mux2_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29404_ _09676_ registers\[21\]\[9\] _13140_ VGND VGND VPWR VPWR _13150_ sky130_fd_sc_hd__mux2_1
XANTENNA_312 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23828_ _09640_ registers\[29\]\[60\] _10016_ VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__mux2_1
XANTENNA_323 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26616_ _11620_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_334 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27596_ registers\[34\]\[15\] _10336_ _12162_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__mux2_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_356 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26547_ _10862_ registers\[42\]\[63\] _11513_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__mux2_1
X_29335_ _09775_ registers\[22\]\[40\] _13113_ VGND VGND VPWR VPWR _13114_ sky130_fd_sc_hd__mux2_1
XANTENNA_367 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_378 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23759_ _09571_ registers\[29\]\[27\] _10039_ VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__mux2_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_389 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16300_ _14592_ VGND VGND VPWR VPWR _14808_ sky130_fd_sc_hd__buf_6
XFILLER_14_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17280_ _15755_ _15759_ _15620_ _15621_ VGND VGND VPWR VPWR _15760_ sky130_fd_sc_hd__o211a_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29266_ _13077_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__clkbuf_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26478_ _11513_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__buf_4
XFILLER_202_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16231_ registers\[24\]\[4\] registers\[25\]\[4\] registers\[26\]\[4\] registers\[27\]\[4\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14741_ sky130_fd_sc_hd__mux4_1
X_28217_ _12494_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__clkbuf_1
X_25429_ _10833_ registers\[50\]\[49\] _10981_ VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__mux2_1
X_29197_ net42 VGND VGND VPWR VPWR _13033_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16162_ _14670_ _14673_ _14585_ VGND VGND VPWR VPWR _14674_ sky130_fd_sc_hd__o21ba_1
XFILLER_166_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28148_ _12458_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__clkbuf_1
X_28079_ _11839_ registers\[31\]\[52\] _12419_ VGND VGND VPWR VPWR _12422_ sky130_fd_sc_hd__mux2_1
X_16093_ _14543_ VGND VGND VPWR VPWR _14607_ sky130_fd_sc_hd__buf_12
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30110_ _13521_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19921_ registers\[44\]\[44\] registers\[45\]\[44\] registers\[46\]\[44\] registers\[47\]\[44\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__mux4_1
X_31090_ _13992_ VGND VGND VPWR VPWR _14037_ sky130_fd_sc_hd__buf_4
XFILLER_170_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30041_ registers\[17\]\[55\] _13050_ _13479_ VGND VGND VPWR VPWR _13485_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19852_ registers\[32\]\[42\] registers\[33\]\[42\] registers\[34\]\[42\] registers\[35\]\[42\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_150_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_150_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18803_ registers\[48\]\[12\] registers\[49\]\[12\] registers\[50\]\[12\] registers\[51\]\[12\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__mux4_1
XFILLER_116_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19783_ registers\[56\]\[40\] registers\[57\]\[40\] registers\[58\]\[40\] registers\[59\]\[40\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__mux4_1
X_16995_ registers\[8\]\[26\] registers\[9\]\[26\] registers\[10\]\[26\] registers\[11\]\[26\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15483_ sky130_fd_sc_hd__mux4_1
X_33800_ clknet_leaf_243_CLK _01914_ VGND VGND VPWR VPWR registers\[40\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18734_ _05111_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__buf_6
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34780_ clknet_leaf_5_CLK _02894_ VGND VGND VPWR VPWR registers\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31992_ clknet_leaf_23_CLK _00164_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
XTAP_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33731_ clknet_leaf_249_CLK _01845_ VGND VGND VPWR VPWR registers\[41\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18665_ registers\[0\]\[8\] registers\[1\]\[8\] registers\[2\]\[8\] registers\[3\]\[8\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__mux4_1
X_30943_ registers\[10\]\[34\] _13006_ _13955_ VGND VGND VPWR VPWR _13960_ sky130_fd_sc_hd__mux2_1
XFILLER_224_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _04376_ _04383_ _04392_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or4_2
X_33662_ clknet_leaf_273_CLK _01776_ VGND VGND VPWR VPWR registers\[42\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30874_ registers\[10\]\[1\] _12937_ _13922_ VGND VGND VPWR VPWR _13924_ sky130_fd_sc_hd__mux2_1
X_18596_ _05130_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__buf_4
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35401_ clknet_leaf_156_CLK _03515_ VGND VGND VPWR VPWR registers\[15\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32613_ clknet_leaf_441_CLK _00727_ VGND VGND VPWR VPWR registers\[58\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17547_ _04332_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_233_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33593_ clknet_leaf_280_CLK _01707_ VGND VGND VPWR VPWR registers\[43\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_890 _09628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35332_ clknet_leaf_223_CLK _03446_ VGND VGND VPWR VPWR registers\[16\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32544_ clknet_leaf_473_CLK _00658_ VGND VGND VPWR VPWR registers\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_17478_ registers\[44\]\[40\] registers\[45\]\[40\] registers\[46\]\[40\] registers\[47\]\[40\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _15952_ sky130_fd_sc_hd__mux4_1
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19217_ _05890_ _05954_ _05955_ _05893_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__a22o_1
X_35263_ clknet_leaf_189_CLK _03377_ VGND VGND VPWR VPWR registers\[17\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_16429_ _14863_ _14931_ _14932_ _14867_ VGND VGND VPWR VPWR _14933_ sky130_fd_sc_hd__a22o_1
XFILLER_177_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32475_ clknet_leaf_58_CLK _00589_ VGND VGND VPWR VPWR registers\[60\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34214_ clknet_leaf_432_CLK _02328_ VGND VGND VPWR VPWR registers\[33\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31426_ _09672_ registers\[6\]\[7\] _14206_ VGND VGND VPWR VPWR _14214_ sky130_fd_sc_hd__mux2_1
X_19148_ _05883_ _05886_ _05887_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__a22o_1
X_35194_ clknet_leaf_185_CLK _03308_ VGND VGND VPWR VPWR registers\[18\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34145_ clknet_leaf_41_CLK _02259_ VGND VGND VPWR VPWR registers\[34\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31357_ _14177_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__clkbuf_1
X_19079_ _05747_ _05820_ _05821_ _05753_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__a22o_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21110_ registers\[0\]\[12\] registers\[1\]\[12\] registers\[2\]\[12\] registers\[3\]\[12\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__mux4_1
X_30308_ _13625_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22090_ _07340_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__clkbuf_4
X_34076_ clknet_leaf_23_CLK _02190_ VGND VGND VPWR VPWR registers\[35\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_31288_ _14141_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33027_ clknet_leaf_269_CLK _01141_ VGND VGND VPWR VPWR registers\[52\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21041_ _07369_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_141_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_141_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30239_ _13589_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24800_ _09594_ registers\[54\]\[38\] _10620_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__mux2_1
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25780_ _10770_ registers\[47\]\[19\] _11170_ VGND VGND VPWR VPWR _11180_ sky130_fd_sc_hd__mux2_1
XFILLER_189_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34978_ clknet_leaf_471_CLK _03092_ VGND VGND VPWR VPWR registers\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_22992_ _09590_ registers\[62\]\[36\] _09578_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__mux2_1
XFILLER_67_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24731_ _09525_ registers\[54\]\[5\] _10587_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__mux2_1
X_33929_ clknet_leaf_236_CLK _02043_ VGND VGND VPWR VPWR registers\[38\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21943_ _07333_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__buf_4
XFILLER_83_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27450_ _12090_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24662_ _10555_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21874_ registers\[48\]\[34\] registers\[49\]\[34\] registers\[50\]\[34\] registers\[51\]\[34\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__mux4_1
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26401_ _11506_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ registers\[61\]\[23\] _09730_ _09965_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__mux2_1
X_20825_ registers\[12\]\[4\] registers\[13\]\[4\] registers\[14\]\[4\] registers\[15\]\[4\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__mux4_1
X_27381_ registers\[36\]\[42\] _10393_ _12051_ VGND VGND VPWR VPWR _12054_ sky130_fd_sc_hd__mux2_1
XFILLER_196_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24593_ _10519_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26332_ _11470_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_1
X_29120_ net15 VGND VGND VPWR VPWR _12981_ sky130_fd_sc_hd__buf_2
X_23544_ _09931_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
X_20756_ registers\[8\]\[2\] registers\[9\]\[2\] registers\[10\]\[2\] registers\[11\]\[2\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__mux4_1
XFILLER_211_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29051_ _09656_ _12933_ VGND VGND VPWR VPWR _12934_ sky130_fd_sc_hd__nor2_8
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26263_ _10848_ registers\[44\]\[56\] _11427_ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__mux2_1
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23475_ _09895_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20687_ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__buf_4
X_25214_ _10754_ registers\[51\]\[11\] _10876_ VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__mux2_1
X_28002_ _12381_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22426_ registers\[40\]\[50\] registers\[41\]\[50\] registers\[42\]\[50\] registers\[43\]\[50\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__mux4_1
X_26194_ _10779_ registers\[44\]\[23\] _11394_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__mux2_1
XFILLER_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25145_ _10834_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22357_ registers\[44\]\[48\] registers\[45\]\[48\] registers\[46\]\[48\] registers\[47\]\[48\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__mux4_1
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_380_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_380_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21308_ _07285_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29953_ registers\[17\]\[13\] _12962_ _13435_ VGND VGND VPWR VPWR _13439_ sky130_fd_sc_hd__mux2_1
X_25076_ _10787_ registers\[52\]\[27\] _10773_ VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__mux2_1
X_22288_ registers\[36\]\[46\] registers\[37\]\[46\] registers\[38\]\[46\] registers\[39\]\[46\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__mux4_1
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28904_ _12855_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24027_ _09567_ registers\[5\]\[25\] _10183_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_132_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_132_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21239_ _07648_ _07918_ _07921_ _07652_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__a22o_1
XFILLER_137_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29884_ _13402_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28835_ _12819_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28766_ _11851_ registers\[26\]\[58\] _12774_ VGND VGND VPWR VPWR _12783_ sky130_fd_sc_hd__mux2_1
XFILLER_120_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16780_ registers\[60\]\[20\] registers\[61\]\[20\] registers\[62\]\[20\] registers\[63\]\[20\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15274_ sky130_fd_sc_hd__mux4_1
X_25978_ _10833_ registers\[46\]\[49\] _11274_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__mux2_1
XFILLER_24_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27717_ _12231_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__clkbuf_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24929_ _09588_ registers\[53\]\[35\] _10691_ VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__mux2_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28697_ _11782_ registers\[26\]\[25\] _12741_ VGND VGND VPWR VPWR _12747_ sky130_fd_sc_hd__mux2_1
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ registers\[48\]\[2\] registers\[49\]\[2\] registers\[50\]\[2\] registers\[51\]\[2\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__mux4_1
XFILLER_98_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27648_ _12150_ VGND VGND VPWR VPWR _12195_ sky130_fd_sc_hd__buf_4
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_131 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_142 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ registers\[40\]\[38\] registers\[41\]\[38\] registers\[42\]\[38\] registers\[43\]\[38\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15877_ sky130_fd_sc_hd__mux4_1
XANTENNA_153 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_199_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_199_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18381_ _05143_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__buf_4
XANTENNA_164 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27579_ registers\[34\]\[7\] _10319_ _12151_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__mux2_1
XANTENNA_175 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_186 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29318_ _09758_ registers\[22\]\[32\] _13102_ VGND VGND VPWR VPWR _13105_ sky130_fd_sc_hd__mux2_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ registers\[32\]\[36\] registers\[33\]\[36\] registers\[34\]\[36\] registers\[35\]\[36\]
+ _15574_ _15575_ VGND VGND VPWR VPWR _15810_ sky130_fd_sc_hd__mux4_1
X_30590_ _09817_ registers\[13\]\[59\] _13764_ VGND VGND VPWR VPWR _13774_ sky130_fd_sc_hd__mux2_1
XFILLER_198_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29249_ _09866_ _10585_ VGND VGND VPWR VPWR _13068_ sky130_fd_sc_hd__nand2_8
X_17263_ _15720_ _15727_ _15736_ _15743_ VGND VGND VPWR VPWR _15744_ sky130_fd_sc_hd__or4_4
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19002_ _05076_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__clkbuf_4
X_16214_ registers\[56\]\[4\] registers\[57\]\[4\] registers\[58\]\[4\] registers\[59\]\[4\]
+ _14723_ _14532_ VGND VGND VPWR VPWR _14724_ sky130_fd_sc_hd__mux4_1
X_32260_ clknet_leaf_253_CLK _00374_ VGND VGND VPWR VPWR registers\[39\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_17194_ _15676_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16145_ registers\[36\]\[2\] registers\[37\]\[2\] registers\[38\]\[2\] registers\[39\]\[2\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14657_ sky130_fd_sc_hd__mux4_1
XFILLER_128_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31211_ registers\[8\]\[33\] net27 _14097_ VGND VGND VPWR VPWR _14101_ sky130_fd_sc_hd__mux2_1
X_32191_ clknet_leaf_460_CLK _00305_ VGND VGND VPWR VPWR registers\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_371_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_371_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16076_ _14578_ VGND VGND VPWR VPWR _14590_ sky130_fd_sc_hd__buf_4
X_31142_ registers\[8\]\[0\] net1 _14064_ VGND VGND VPWR VPWR _14065_ sky130_fd_sc_hd__mux2_1
XFILLER_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19904_ _05069_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__buf_4
X_31073_ _14028_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__clkbuf_1
X_35950_ clknet_leaf_391_CLK _04064_ VGND VGND VPWR VPWR registers\[6\]\[32\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_123_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_123_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_30__f_CLK clknet_5_15_0_CLK VGND VGND VPWR VPWR clknet_6_30__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34901_ clknet_leaf_97_CLK _03015_ VGND VGND VPWR VPWR registers\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_30024_ registers\[17\]\[47\] _13033_ _13468_ VGND VGND VPWR VPWR _13476_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19835_ registers\[12\]\[41\] registers\[13\]\[41\] registers\[14\]\[41\] registers\[15\]\[41\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__mux4_1
X_35881_ clknet_leaf_400_CLK _03995_ VGND VGND VPWR VPWR registers\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34832_ clknet_leaf_115_CLK _02946_ VGND VGND VPWR VPWR registers\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19766_ _06182_ _06488_ _06489_ _06185_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__a22o_1
X_16978_ registers\[40\]\[26\] registers\[41\]\[26\] registers\[42\]\[26\] registers\[43\]\[26\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15466_ sky130_fd_sc_hd__mux4_1
XFILLER_77_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 DW[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_8
XFILLER_65_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18717_ _05051_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__buf_4
X_34763_ clknet_leaf_152_CLK _02877_ VGND VGND VPWR VPWR registers\[25\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19697_ _06187_ _06421_ _06422_ _06192_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__a22o_1
X_31975_ clknet_leaf_6_CLK _00145_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
X_33714_ clknet_leaf_360_CLK _01828_ VGND VGND VPWR VPWR registers\[41\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_18648_ _05399_ _05402_ _05074_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__o21ba_2
X_30926_ registers\[10\]\[26\] _12989_ _13944_ VGND VGND VPWR VPWR _13951_ sky130_fd_sc_hd__mux2_1
X_34694_ clknet_leaf_218_CLK _02808_ VGND VGND VPWR VPWR registers\[26\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33645_ clknet_leaf_330_CLK _01759_ VGND VGND VPWR VPWR registers\[42\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_30857_ _13914_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__clkbuf_1
X_18579_ registers\[56\]\[6\] registers\[57\]\[6\] registers\[58\]\[6\] registers\[59\]\[6\]
+ _05272_ _05081_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__mux4_1
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20610_ net75 net76 VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__or2b_4
X_33576_ clknet_leaf_430_CLK _01690_ VGND VGND VPWR VPWR registers\[43\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_21590_ _07333_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__buf_6
X_30788_ _13878_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35315_ clknet_leaf_409_CLK _03429_ VGND VGND VPWR VPWR registers\[16\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_20541_ _05119_ _07240_ _07241_ _05131_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__a22o_1
X_32527_ clknet_leaf_139_CLK _00641_ VGND VGND VPWR VPWR registers\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35246_ clknet_leaf_397_CLK _03360_ VGND VGND VPWR VPWR registers\[17\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_23260_ _09768_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
X_20472_ registers\[12\]\[60\] registers\[13\]\[60\] registers\[14\]\[60\] registers\[15\]\[60\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__mux4_1
X_32458_ clknet_leaf_165_CLK _00572_ VGND VGND VPWR VPWR registers\[29\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22211_ _08761_ _08865_ _08866_ _08764_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__a22o_1
X_31409_ _14204_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__clkbuf_1
X_35177_ clknet_leaf_404_CLK _03291_ VGND VGND VPWR VPWR registers\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_362_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_362_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23191_ registers\[9\]\[13\] _09685_ _09722_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__mux2_1
X_32389_ clknet_leaf_202_CLK _00503_ VGND VGND VPWR VPWR registers\[61\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34128_ clknet_leaf_128_CLK _02242_ VGND VGND VPWR VPWR registers\[34\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_22142_ registers\[28\]\[41\] registers\[29\]\[41\] registers\[30\]\[41\] registers\[31\]\[41\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34059_ clknet_leaf_165_CLK _02173_ VGND VGND VPWR VPWR registers\[36\]\[61\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_114_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_114_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22073_ registers\[40\]\[40\] registers\[41\]\[40\] registers\[42\]\[40\] registers\[43\]\[40\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__mux4_1
X_26950_ net36 VGND VGND VPWR VPWR _11816_ sky130_fd_sc_hd__clkbuf_4
XTAP_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21024_ registers\[56\]\[10\] registers\[57\]\[10\] registers\[58\]\[10\] registers\[59\]\[10\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__mux4_1
X_25901_ _10756_ registers\[46\]\[12\] _11241_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__mux2_1
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26881_ net11 VGND VGND VPWR VPWR _11769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28620_ _12706_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25832_ _11207_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28551_ _12647_ VGND VGND VPWR VPWR _12670_ sky130_fd_sc_hd__buf_4
X_25763_ _11171_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
X_22975_ _09579_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
X_27502_ _12117_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__clkbuf_1
X_24714_ _10582_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
X_21926_ registers\[20\]\[35\] registers\[21\]\[35\] registers\[22\]\[35\] registers\[23\]\[35\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__mux4_1
XFILLER_216_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28482_ _11837_ registers\[28\]\[51\] _12632_ VGND VGND VPWR VPWR _12634_ sky130_fd_sc_hd__mux2_1
X_25694_ registers\[48\]\[43\] _10395_ _11130_ VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__mux2_1
XFILLER_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27433_ _12081_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__clkbuf_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24645_ _10546_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ registers\[16\]\[33\] registers\[17\]\[33\] registers\[18\]\[33\] registers\[19\]\[33\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__mux4_1
XFILLER_43_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20808_ _07433_ _07501_ _07502_ _07438_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__a22o_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24576_ _10508_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
X_27364_ registers\[36\]\[34\] _10376_ _12040_ VGND VGND VPWR VPWR _12045_ sky130_fd_sc_hd__mux2_1
X_21788_ _08418_ _08454_ _08455_ _08421_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__a22o_1
XFILLER_243_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29103_ _12969_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23527_ _09922_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26315_ _11461_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
X_20739_ registers\[40\]\[2\] registers\[41\]\[2\] registers\[42\]\[2\] registers\[43\]\[2\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__mux4_1
X_27295_ registers\[36\]\[1\] _10307_ _12007_ VGND VGND VPWR VPWR _12009_ sky130_fd_sc_hd__mux2_1
XFILLER_211_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29034_ registers\[24\]\[57\] _10424_ _12916_ VGND VGND VPWR VPWR _12924_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26246_ _10831_ registers\[44\]\[48\] _11416_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__mux2_1
XFILLER_167_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23458_ _09886_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22409_ _09055_ _09058_ _08748_ _08749_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__o211a_1
X_26177_ _10762_ registers\[44\]\[15\] _11383_ VGND VGND VPWR VPWR _11389_ sky130_fd_sc_hd__mux2_1
XFILLER_104_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23389_ _09848_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_353_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_353_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25128_ net39 VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__buf_2
XFILLER_178_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29936_ registers\[17\]\[5\] _12945_ _13424_ VGND VGND VPWR VPWR _13430_ sky130_fd_sc_hd__mux2_1
X_17950_ registers\[52\]\[53\] registers\[53\]\[53\] registers\[54\]\[53\] registers\[55\]\[53\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_105_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_105_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ _10776_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_991 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16901_ _15144_ _15390_ _15391_ _15147_ VGND VGND VPWR VPWR _15392_ sky130_fd_sc_hd__a22o_1
XFILLER_78_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17881_ registers\[60\]\[51\] registers\[61\]\[51\] registers\[62\]\[51\] registers\[63\]\[51\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__mux4_1
X_29867_ _13393_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19620_ _06036_ _06346_ _06347_ _06039_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__a22o_1
X_16832_ _15321_ _15324_ _15288_ VGND VGND VPWR VPWR _15325_ sky130_fd_sc_hd__o21ba_1
X_28818_ _12810_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29798_ _13357_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19551_ _05069_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__buf_4
X_28749_ _12718_ VGND VGND VPWR VPWR _12774_ sky130_fd_sc_hd__buf_4
X_16763_ _14952_ _15256_ _15257_ _14957_ VGND VGND VPWR VPWR _15258_ sky130_fd_sc_hd__a22o_1
XFILLER_219_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18502_ _05150_ _05260_ _05261_ _05160_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__a22o_1
XFILLER_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19482_ registers\[12\]\[31\] registers\[13\]\[31\] registers\[14\]\[31\] registers\[15\]\[31\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__mux4_1
X_31760_ _14389_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16694_ _15190_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30711_ registers\[12\]\[52\] _13044_ _13835_ VGND VGND VPWR VPWR _13838_ sky130_fd_sc_hd__mux2_1
X_18433_ _05191_ _05194_ _05163_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31691_ _14353_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__clkbuf_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33430_ clknet_leaf_123_CLK _01544_ VGND VGND VPWR VPWR registers\[45\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30642_ _13801_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__clkbuf_1
X_18364_ _05080_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ registers\[8\]\[35\] registers\[9\]\[35\] registers\[10\]\[35\] registers\[11\]\[35\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15794_ sky130_fd_sc_hd__mux4_1
XFILLER_72_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33361_ clknet_leaf_129_CLK _01475_ VGND VGND VPWR VPWR registers\[46\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30573_ _13765_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__clkbuf_1
X_18295_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__buf_2
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35100_ clknet_leaf_478_CLK _03214_ VGND VGND VPWR VPWR registers\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32312_ clknet_leaf_428_CLK _00426_ VGND VGND VPWR VPWR registers\[19\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17246_ _15723_ _15726_ _15620_ _15621_ VGND VGND VPWR VPWR _15727_ sky130_fd_sc_hd__o211a_1
X_36080_ clknet_leaf_366_CLK _04194_ VGND VGND VPWR VPWR registers\[59\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_33292_ clknet_leaf_168_CLK _01406_ VGND VGND VPWR VPWR registers\[48\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35031_ clknet_leaf_103_CLK _03145_ VGND VGND VPWR VPWR registers\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_32243_ clknet_leaf_348_CLK _00357_ VGND VGND VPWR VPWR registers\[39\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17177_ _15549_ _15658_ _15659_ _15553_ VGND VGND VPWR VPWR _15660_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_344_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_344_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16128_ registers\[16\]\[1\] registers\[17\]\[1\] registers\[18\]\[1\] registers\[19\]\[1\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14641_ sky130_fd_sc_hd__mux4_1
XFILLER_227_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32174_ clknet_leaf_86_CLK _00288_ VGND VGND VPWR VPWR registers\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31125_ _14055_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16059_ _14495_ VGND VGND VPWR VPWR _14573_ sky130_fd_sc_hd__buf_12
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31056_ _14019_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__clkbuf_1
X_35933_ clknet_leaf_476_CLK _04047_ VGND VGND VPWR VPWR registers\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30007_ registers\[17\]\[39\] _13016_ _13457_ VGND VGND VPWR VPWR _13467_ sky130_fd_sc_hd__mux2_1
X_19818_ registers\[40\]\[41\] registers\[41\]\[41\] registers\[42\]\[41\] registers\[43\]\[41\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__mux4_1
XFILLER_233_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35864_ clknet_leaf_474_CLK _03978_ VGND VGND VPWR VPWR registers\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34815_ clknet_leaf_197_CLK _02929_ VGND VGND VPWR VPWR registers\[24\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_19749_ _06469_ _06472_ _06161_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__o21ba_1
X_35795_ clknet_leaf_79_CLK _03909_ VGND VGND VPWR VPWR registers\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_22760_ _09155_ _09397_ _09398_ _09158_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__a22o_1
X_34746_ clknet_leaf_184_CLK _02860_ VGND VGND VPWR VPWR registers\[25\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31958_ clknet_leaf_0_CLK _00190_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21711_ registers\[24\]\[29\] registers\[25\]\[29\] registers\[26\]\[29\] registers\[27\]\[29\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__mux4_1
X_30909_ registers\[10\]\[18\] _12972_ _13933_ VGND VGND VPWR VPWR _13942_ sky130_fd_sc_hd__mux2_1
X_22691_ _09109_ _09331_ _09332_ _09114_ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__a22o_1
X_34677_ clknet_leaf_413_CLK _02791_ VGND VGND VPWR VPWR registers\[26\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31889_ _14457_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__clkbuf_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24430_ _10429_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21642_ registers\[28\]\[27\] registers\[29\]\[27\] registers\[30\]\[27\] registers\[31\]\[27\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__mux4_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33628_ clknet_leaf_27_CLK _01742_ VGND VGND VPWR VPWR registers\[42\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24361_ registers\[57\]\[37\] _10382_ _10368_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__mux2_1
X_33559_ clknet_leaf_128_CLK _01673_ VGND VGND VPWR VPWR registers\[43\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ registers\[20\]\[25\] registers\[21\]\[25\] registers\[22\]\[25\] registers\[23\]\[25\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__mux4_1
XANTENNA_31 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26100_ _11348_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
X_23312_ _09803_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_42 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20524_ _05136_ _07223_ _07224_ _05146_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__a22o_1
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_53 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27080_ _11895_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_64 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24292_ net7 VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__buf_4
XANTENNA_75 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26031_ _11300_ VGND VGND VPWR VPWR _11312_ sky130_fd_sc_hd__buf_4
XANTENNA_86 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23243_ _09757_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
X_35229_ clknet_leaf_5_CLK _03343_ VGND VGND VPWR VPWR registers\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_20455_ registers\[40\]\[60\] registers\[41\]\[60\] registers\[42\]\[60\] registers\[43\]\[60\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__mux4_1
XFILLER_197_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_335_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_335_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23174_ _09716_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20386_ registers\[24\]\[57\] registers\[25\]\[57\] registers\[26\]\[57\] registers\[27\]\[57\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__mux4_1
XFILLER_107_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22125_ registers\[56\]\[41\] registers\[57\]\[41\] registers\[58\]\[41\] registers\[59\]\[41\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__mux4_1
XTAP_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27982_ _11742_ registers\[31\]\[6\] _12364_ VGND VGND VPWR VPWR _12371_ sky130_fd_sc_hd__mux2_1
Xoutput160 net160 VGND VGND VPWR VPWR D2[15] sky130_fd_sc_hd__buf_2
XTAP_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput171 net171 VGND VGND VPWR VPWR D2[25] sky130_fd_sc_hd__buf_2
XFILLER_82_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput182 net182 VGND VGND VPWR VPWR D2[35] sky130_fd_sc_hd__buf_2
X_29721_ registers\[1\]\[31\] _13000_ _13315_ VGND VGND VPWR VPWR _13317_ sky130_fd_sc_hd__mux2_1
XTAP_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput193 net193 VGND VGND VPWR VPWR D2[45] sky130_fd_sc_hd__buf_2
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26933_ _11804_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__clkbuf_1
X_22056_ _08712_ _08715_ _08405_ _08406_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__o211a_1
XTAP_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21007_ _07373_ _07695_ _07696_ _07383_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__a22o_1
XFILLER_88_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29652_ registers\[20\]\[63\] _13066_ _13210_ VGND VGND VPWR VPWR _13280_ sky130_fd_sc_hd__mux2_1
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26864_ _11757_ registers\[3\]\[13\] _11751_ VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_236_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28603_ _12697_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25815_ _11198_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29583_ _13210_ VGND VGND VPWR VPWR _13244_ sky130_fd_sc_hd__buf_4
XFILLER_60_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26795_ registers\[40\]\[51\] _10412_ _11713_ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__mux2_1
X_28534_ _12661_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__clkbuf_1
X_25746_ _11162_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22958_ _09567_ registers\[62\]\[25\] _09557_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__mux2_1
XFILLER_90_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21909_ registers\[60\]\[35\] registers\[61\]\[35\] registers\[62\]\[35\] registers\[63\]\[35\]
+ _08541_ _08335_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__mux4_1
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28465_ _11820_ registers\[28\]\[43\] _12621_ VGND VGND VPWR VPWR _12625_ sky130_fd_sc_hd__mux2_1
XFILLER_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22889_ net34 VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__clkbuf_4
X_25677_ registers\[48\]\[35\] _10378_ _11119_ VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__mux2_1
XFILLER_203_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27416_ registers\[36\]\[59\] _10428_ _12062_ VGND VGND VPWR VPWR _12072_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24628_ _09559_ registers\[55\]\[21\] _10536_ VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__mux2_1
XFILLER_203_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28396_ _11750_ registers\[28\]\[10\] _12588_ VGND VGND VPWR VPWR _12589_ sky130_fd_sc_hd__mux2_1
XFILLER_197_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24559_ _09628_ registers\[56\]\[54\] _10495_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__mux2_1
XFILLER_200_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27347_ registers\[36\]\[26\] _10359_ _12029_ VGND VGND VPWR VPWR _12036_ sky130_fd_sc_hd__mux2_1
XFILLER_223_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17100_ registers\[60\]\[29\] registers\[61\]\[29\] registers\[62\]\[29\] registers\[63\]\[29\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15585_ sky130_fd_sc_hd__mux4_1
X_18080_ registers\[0\]\[57\] registers\[1\]\[57\] registers\[2\]\[57\] registers\[3\]\[57\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__mux4_1
X_27278_ _11999_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29017_ registers\[24\]\[49\] _10407_ _12905_ VGND VGND VPWR VPWR _12915_ sky130_fd_sc_hd__mux2_1
X_17031_ _15514_ _15517_ _15277_ _15278_ VGND VGND VPWR VPWR _15518_ sky130_fd_sc_hd__o211a_1
X_26229_ _11371_ VGND VGND VPWR VPWR _11416_ sky130_fd_sc_hd__buf_4
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_326_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_326_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18982_ registers\[12\]\[17\] registers\[13\]\[17\] registers\[14\]\[17\] registers\[15\]\[17\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__mux4_1
XFILLER_139_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29919_ _13420_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__clkbuf_1
X_17933_ registers\[28\]\[52\] registers\[29\]\[52\] registers\[30\]\[52\] registers\[31\]\[52\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__mux4_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32930_ clknet_leaf_443_CLK _01044_ VGND VGND VPWR VPWR registers\[53\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17864_ registers\[20\]\[50\] registers\[21\]\[50\] registers\[22\]\[50\] registers\[23\]\[50\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__mux4_1
XFILLER_152_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19603_ registers\[36\]\[35\] registers\[37\]\[35\] registers\[38\]\[35\] registers\[39\]\[35\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__mux4_1
XFILLER_113_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16815_ registers\[44\]\[21\] registers\[45\]\[21\] registers\[46\]\[21\] registers\[47\]\[21\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15308_ sky130_fd_sc_hd__mux4_1
XFILLER_187_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32861_ clknet_leaf_55_CLK _00975_ VGND VGND VPWR VPWR registers\[54\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17795_ _14502_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__clkbuf_8
XFILLER_47_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34600_ clknet_leaf_453_CLK _02714_ VGND VGND VPWR VPWR registers\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31812_ _14416_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__clkbuf_1
X_19534_ registers\[32\]\[33\] registers\[33\]\[33\] registers\[34\]\[33\] registers\[35\]\[33\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__mux4_1
X_35580_ clknet_leaf_299_CLK _03694_ VGND VGND VPWR VPWR registers\[12\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_16746_ _15198_ _15239_ _15240_ _15204_ VGND VGND VPWR VPWR _15241_ sky130_fd_sc_hd__a22o_1
X_32792_ clknet_leaf_67_CLK _00906_ VGND VGND VPWR VPWR registers\[55\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34531_ clknet_leaf_473_CLK _02645_ VGND VGND VPWR VPWR registers\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31743_ _14380_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__clkbuf_1
X_19465_ registers\[40\]\[31\] registers\[41\]\[31\] registers\[42\]\[31\] registers\[43\]\[31\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__mux4_1
X_16677_ _14863_ _15172_ _15173_ _14867_ VGND VGND VPWR VPWR _15174_ sky130_fd_sc_hd__a22o_1
XFILLER_22_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18416_ registers\[60\]\[1\] registers\[61\]\[1\] registers\[62\]\[1\] registers\[63\]\[1\]
+ _05091_ _05093_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__mux4_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34462_ clknet_leaf_487_CLK _02576_ VGND VGND VPWR VPWR registers\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31674_ registers\[63\]\[61\] net58 _14276_ VGND VGND VPWR VPWR _14344_ sky130_fd_sc_hd__mux2_1
X_19396_ _06126_ _06129_ _05818_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36201_ clknet_leaf_92_CLK _00083_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dfxtp_1
X_33413_ clknet_leaf_256_CLK _01527_ VGND VGND VPWR VPWR registers\[46\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18347_ registers\[8\]\[0\] registers\[9\]\[0\] registers\[10\]\[0\] registers\[11\]\[0\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__mux4_1
X_30625_ registers\[12\]\[11\] _12958_ _13791_ VGND VGND VPWR VPWR _13793_ sky130_fd_sc_hd__mux2_1
XFILLER_226_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34393_ clknet_leaf_21_CLK _02507_ VGND VGND VPWR VPWR registers\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36132_ clknet_leaf_440_CLK _04246_ VGND VGND VPWR VPWR registers\[49\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_33344_ clknet_leaf_257_CLK _01458_ VGND VGND VPWR VPWR registers\[47\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_18278_ net77 VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__buf_6
XFILLER_198_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30556_ _13756_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput40 DW[45] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
X_17229_ _15638_ _15709_ _15710_ _15643_ VGND VGND VPWR VPWR _15711_ sky130_fd_sc_hd__a22o_1
X_36063_ clknet_leaf_42_CLK _04177_ VGND VGND VPWR VPWR registers\[59\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33275_ clknet_leaf_281_CLK _01389_ VGND VGND VPWR VPWR registers\[48\]\[45\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_317_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_317_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30487_ _13708_ VGND VGND VPWR VPWR _13720_ sky130_fd_sc_hd__buf_4
Xinput51 DW[55] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_16
Xinput62 DW[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
Xinput73 R2[2] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
X_35014_ clknet_leaf_208_CLK _03128_ VGND VGND VPWR VPWR registers\[21\]\[56\] sky130_fd_sc_hd__dfxtp_1
Xinput84 RW[1] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_6
X_20240_ registers\[32\]\[53\] registers\[33\]\[53\] registers\[34\]\[53\] registers\[35\]\[53\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__mux4_1
X_32226_ clknet_leaf_424_CLK _00340_ VGND VGND VPWR VPWR registers\[39\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20171_ registers\[40\]\[51\] registers\[41\]\[51\] registers\[42\]\[51\] registers\[43\]\[51\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__mux4_1
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32157_ clknet_leaf_27_CLK _00271_ VGND VGND VPWR VPWR registers\[39\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31108_ _14046_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32088_ clknet_leaf_489_CLK _00001_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35916_ clknet_leaf_143_CLK _04030_ VGND VGND VPWR VPWR registers\[7\]\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23930_ _10137_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
X_31039_ _14010_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ _10101_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35847_ clknet_leaf_216_CLK _03961_ VGND VGND VPWR VPWR registers\[8\]\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25600_ net85 net84 _10584_ VGND VGND VPWR VPWR _11083_ sky130_fd_sc_hd__or3_1
X_22812_ _09446_ _09449_ _07398_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__o21ba_1
XFILLER_244_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23792_ _10064_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_708 _07295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26580_ _11601_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__clkbuf_1
X_35778_ clknet_leaf_241_CLK _03892_ VGND VGND VPWR VPWR registers\[0\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_719 _07338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22743_ registers\[4\]\[59\] registers\[5\]\[59\] registers\[6\]\[59\] registers\[7\]\[59\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25531_ registers\[4\]\[31\] _10370_ _11045_ VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__mux2_1
X_34729_ clknet_leaf_406_CLK _02843_ VGND VGND VPWR VPWR registers\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25462_ _09941_ _10584_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__or2_1
X_28250_ registers\[2\]\[5\] _10315_ _12506_ VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22674_ _09012_ _09314_ _09315_ _09018_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__a22o_1
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24413_ net50 VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__buf_4
XFILLER_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27201_ _11959_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__clkbuf_1
X_21625_ registers\[56\]\[27\] registers\[57\]\[27\] registers\[58\]\[27\] registers\[59\]\[27\]
+ _08194_ _07984_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__mux4_1
XFILLER_244_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25393_ _10972_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__clkbuf_1
X_28181_ _12475_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27132_ _11839_ registers\[38\]\[52\] _11920_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__mux2_1
XFILLER_194_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24344_ _10371_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21556_ registers\[60\]\[25\] registers\[61\]\[25\] registers\[62\]\[25\] registers\[63\]\[25\]
+ _08198_ _07992_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__mux4_1
XFILLER_21_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20507_ registers\[16\]\[61\] registers\[17\]\[61\] registers\[18\]\[61\] registers\[19\]\[61\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__mux4_1
X_27063_ _11886_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24275_ _10324_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_308_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_308_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21487_ registers\[56\]\[23\] registers\[57\]\[23\] registers\[58\]\[23\] registers\[59\]\[23\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__mux4_1
X_26014_ _11303_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
X_23226_ registers\[39\]\[24\] _09740_ _09700_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__mux2_1
X_20438_ _07138_ _07141_ _06855_ _06856_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__o211a_1
XFILLER_181_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23157_ net85 net84 _09654_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__or3_1
XFILLER_136_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20369_ registers\[36\]\[57\] registers\[37\]\[57\] registers\[38\]\[57\] registers\[39\]\[57\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__mux4_1
XFILLER_175_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1107 _14553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22108_ registers\[28\]\[40\] registers\[29\]\[40\] registers\[30\]\[40\] registers\[31\]\[40\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__mux4_1
XTAP_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1118 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23088_ registers\[39\]\[0\] _09648_ _09658_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__mux2_1
XTAP_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27965_ _12361_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1129 _14600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29704_ registers\[1\]\[23\] _12983_ _13304_ VGND VGND VPWR VPWR _13308_ sky130_fd_sc_hd__mux2_1
XFILLER_88_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26916_ _11729_ VGND VGND VPWR VPWR _11793_ sky130_fd_sc_hd__buf_4
X_22039_ _08668_ _08683_ _08692_ _08699_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__or4_1
XTAP_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27896_ _12325_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29635_ _13271_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__clkbuf_1
XTAP_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26847_ net63 VGND VGND VPWR VPWR _11746_ sky130_fd_sc_hd__clkbuf_4
XTAP_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16600_ registers\[56\]\[15\] registers\[57\]\[15\] registers\[58\]\[15\] registers\[59\]\[15\]
+ _15066_ _14856_ VGND VGND VPWR VPWR _15099_ sky130_fd_sc_hd__mux4_1
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17580_ registers\[28\]\[42\] registers\[29\]\[42\] registers\[30\]\[42\] registers\[31\]\[42\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__mux4_1
X_29566_ _13235_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__clkbuf_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26778_ registers\[40\]\[43\] _10395_ _11702_ VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28517_ _12652_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__clkbuf_1
X_16531_ registers\[36\]\[13\] registers\[37\]\[13\] registers\[38\]\[13\] registers\[39\]\[13\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _15032_ sky130_fd_sc_hd__mux4_1
X_25729_ registers\[48\]\[60\] _10430_ _11085_ VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29497_ _09804_ registers\[21\]\[53\] _13195_ VGND VGND VPWR VPWR _13199_ sky130_fd_sc_hd__mux2_1
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19250_ registers\[36\]\[25\] registers\[37\]\[25\] registers\[38\]\[25\] registers\[39\]\[25\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__mux4_1
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16462_ registers\[44\]\[11\] registers\[45\]\[11\] registers\[46\]\[11\] registers\[47\]\[11\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _14965_ sky130_fd_sc_hd__mux4_1
XFILLER_31_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28448_ _11803_ registers\[28\]\[35\] _12610_ VGND VGND VPWR VPWR _12616_ sky130_fd_sc_hd__mux2_1
XFILLER_177_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18201_ _14491_ _04965_ _04966_ _14501_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a22o_1
XFILLER_223_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19181_ registers\[32\]\[23\] registers\[33\]\[23\] registers\[34\]\[23\] registers\[35\]\[23\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__mux4_1
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28379_ _11734_ registers\[28\]\[2\] _12577_ VGND VGND VPWR VPWR _12580_ sky130_fd_sc_hd__mux2_1
X_16393_ _14855_ _14896_ _14897_ _14861_ VGND VGND VPWR VPWR _14898_ sky130_fd_sc_hd__a22o_1
XFILLER_31_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18132_ registers\[56\]\[59\] registers\[57\]\[59\] registers\[58\]\[59\] registers\[59\]\[59\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__mux4_1
XFILLER_19_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30410_ _13679_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31390_ registers\[7\]\[54\] net50 _14190_ VGND VGND VPWR VPWR _14195_ sky130_fd_sc_hd__mux2_1
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18063_ _04812_ _04819_ _04826_ _04833_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__or4_4
X_30341_ _13643_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ _15472_ _15481_ _15492_ _15501_ VGND VGND VPWR VPWR _15502_ sky130_fd_sc_hd__or4_4
X_33060_ clknet_leaf_440_CLK _01174_ VGND VGND VPWR VPWR registers\[51\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_30272_ _13606_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__clkbuf_1
X_32011_ clknet_leaf_29_CLK _00185_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18965_ _05540_ _05709_ _05710_ _05545_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__a22o_1
XANTENNA_1630 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1641 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17916_ _04540_ _04689_ _04690_ _04546_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__a22o_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1652 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33962_ clknet_leaf_427_CLK _02076_ VGND VGND VPWR VPWR registers\[37\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1663 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18896_ registers\[44\]\[15\] registers\[45\]\[15\] registers\[46\]\[15\] registers\[47\]\[15\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__mux4_1
XTAP_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1674 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1685 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32913_ clknet_leaf_174_CLK _01027_ VGND VGND VPWR VPWR registers\[53\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1696 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35701_ clknet_leaf_324_CLK _03815_ VGND VGND VPWR VPWR registers\[10\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17847_ _14573_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__buf_4
X_33893_ clknet_leaf_433_CLK _02007_ VGND VGND VPWR VPWR registers\[38\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32844_ clknet_leaf_142_CLK _00958_ VGND VGND VPWR VPWR registers\[55\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35632_ clknet_leaf_376_CLK _03746_ VGND VGND VPWR VPWR registers\[11\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_17778_ _04481_ _04555_ _04556_ _04484_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__a22o_1
XFILLER_214_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19517_ _06031_ _06246_ _06247_ _06034_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__a22o_1
X_16729_ registers\[28\]\[18\] registers\[29\]\[18\] registers\[30\]\[18\] registers\[31\]\[18\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15225_ sky130_fd_sc_hd__mux4_1
X_35563_ clknet_leaf_397_CLK _03677_ VGND VGND VPWR VPWR registers\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_32775_ clknet_leaf_262_CLK _00889_ VGND VGND VPWR VPWR registers\[56\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34514_ clknet_leaf_99_CLK _02628_ VGND VGND VPWR VPWR registers\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_19448_ _06176_ _06179_ _06180_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__o21ba_1
X_31726_ registers\[59\]\[21\] net14 _14370_ VGND VGND VPWR VPWR _14372_ sky130_fd_sc_hd__mux2_1
XFILLER_165_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35494_ clknet_leaf_461_CLK _03608_ VGND VGND VPWR VPWR registers\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34445_ clknet_leaf_141_CLK _02559_ VGND VGND VPWR VPWR registers\[30\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_31657_ _14335_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__clkbuf_1
X_19379_ registers\[24\]\[28\] registers\[25\]\[28\] registers\[26\]\[28\] registers\[27\]\[28\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_94_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_94_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21410_ _08055_ _08064_ _08074_ _08088_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__or4_4
XFILLER_241_1366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30608_ registers\[12\]\[3\] _12941_ _13780_ VGND VGND VPWR VPWR _13784_ sky130_fd_sc_hd__mux2_1
X_34376_ clknet_leaf_214_CLK _02490_ VGND VGND VPWR VPWR registers\[31\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22390_ _08766_ _09039_ _09040_ _08771_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__a22o_1
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31588_ _14276_ VGND VGND VPWR VPWR _14299_ sky130_fd_sc_hd__buf_4
XFILLER_148_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36115_ clknet_leaf_70_CLK _04229_ VGND VGND VPWR VPWR registers\[49\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33327_ clknet_leaf_362_CLK _01441_ VGND VGND VPWR VPWR registers\[47\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_21341_ registers\[36\]\[19\] registers\[37\]\[19\] registers\[38\]\[19\] registers\[39\]\[19\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__mux4_1
XFILLER_108_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30539_ _13747_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36046_ clknet_leaf_173_CLK _04160_ VGND VGND VPWR VPWR registers\[59\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_24060_ _10206_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
X_33258_ clknet_leaf_424_CLK _01372_ VGND VGND VPWR VPWR registers\[48\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_21272_ registers\[56\]\[17\] registers\[57\]\[17\] registers\[58\]\[17\] registers\[59\]\[17\]
+ _07851_ _07641_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__mux4_1
XFILLER_191_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23011_ _09603_ registers\[62\]\[42\] _09599_ VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__mux2_1
X_20223_ _06717_ _06932_ _06933_ _06720_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__a22o_1
XFILLER_116_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32209_ clknet_leaf_318_CLK _00323_ VGND VGND VPWR VPWR registers\[9\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33189_ clknet_leaf_456_CLK _01303_ VGND VGND VPWR VPWR registers\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20154_ _06862_ _06865_ _06866_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__o21ba_1
XFILLER_89_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27750_ registers\[33\]\[24\] _10355_ _12244_ VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__mux2_1
X_24962_ _10714_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
X_20085_ registers\[24\]\[48\] registers\[25\]\[48\] registers\[26\]\[48\] registers\[27\]\[48\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__mux4_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26701_ _11665_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_1
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ _10128_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27681_ _12212_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__clkbuf_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24893_ _09552_ registers\[53\]\[18\] _10669_ VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__mux2_1
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29420_ _13158_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__clkbuf_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26632_ _11628_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__clkbuf_1
X_23844_ _10092_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__clkbuf_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_505 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_516 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_226_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_527 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29351_ _09793_ registers\[22\]\[48\] _13113_ VGND VGND VPWR VPWR _13122_ sky130_fd_sc_hd__mux2_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26563_ _11592_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_538 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23775_ _10055_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
X_20987_ registers\[44\]\[9\] registers\[45\]\[9\] registers\[46\]\[9\] registers\[47\]\[9\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__mux4_1
XFILLER_226_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_549 _04440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28302_ _12505_ VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__buf_4
XFILLER_241_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25514_ registers\[4\]\[23\] _10353_ _11034_ VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__mux2_1
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22726_ registers\[32\]\[59\] registers\[33\]\[59\] registers\[34\]\[59\] registers\[35\]\[59\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__mux4_1
XFILLER_159_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29282_ _09689_ registers\[22\]\[15\] _13080_ VGND VGND VPWR VPWR _13086_ sky130_fd_sc_hd__mux2_1
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26494_ _11555_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28233_ _12502_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22657_ registers\[16\]\[56\] registers\[17\]\[56\] registers\[18\]\[56\] registers\[19\]\[56\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__mux4_1
X_25445_ _10999_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_85_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_85_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_199_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21608_ registers\[16\]\[26\] registers\[17\]\[26\] registers\[18\]\[26\] registers\[19\]\[26\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__mux4_1
XFILLER_185_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28164_ _12466_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__clkbuf_1
X_22588_ registers\[0\]\[54\] registers\[1\]\[54\] registers\[2\]\[54\] registers\[3\]\[54\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__mux4_1
X_25376_ _10963_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_975 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27115_ _11822_ registers\[38\]\[44\] _11909_ VGND VGND VPWR VPWR _11914_ sky130_fd_sc_hd__mux2_1
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21539_ _08075_ _08212_ _08213_ _08078_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__a22o_1
X_24327_ registers\[57\]\[26\] _10359_ _10347_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__mux2_1
X_28095_ _11855_ registers\[31\]\[60\] _12363_ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__mux2_1
XFILLER_154_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24258_ net45 VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__buf_4
X_27046_ _11753_ registers\[38\]\[11\] _11876_ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__mux2_1
X_23209_ registers\[9\]\[20\] _09699_ _09735_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__mux2_1
XFILLER_181_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24189_ _10274_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28997_ _12904_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__clkbuf_1
XTAP_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1068 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18750_ _05079_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__buf_4
X_27948_ registers\[32\]\[54\] _10418_ _12348_ VGND VGND VPWR VPWR _12353_ sky130_fd_sc_hd__mux2_1
XTAP_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ registers\[8\]\[46\] registers\[9\]\[46\] registers\[10\]\[46\] registers\[11\]\[46\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__mux4_1
XFILLER_23_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _05435_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
XTAP_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27879_ registers\[32\]\[21\] _10349_ _12315_ VGND VGND VPWR VPWR _12317_ sky130_fd_sc_hd__mux2_1
XTAP_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29618_ _13262_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__clkbuf_1
X_17632_ _15892_ _04413_ _04414_ _15896_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__a22o_1
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30890_ registers\[10\]\[9\] _12953_ _13922_ VGND VGND VPWR VPWR _13932_ sky130_fd_sc_hd__mux2_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17563_ _15884_ _04346_ _04347_ _15890_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__a22o_1
X_29549_ _13226_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19302_ _05130_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16514_ _14801_ _15014_ _15015_ _14804_ VGND VGND VPWR VPWR _15016_ sky130_fd_sc_hd__a22o_1
XFILLER_147_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32560_ clknet_leaf_375_CLK _00674_ VGND VGND VPWR VPWR registers\[5\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17494_ _14573_ VGND VGND VPWR VPWR _15968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31511_ _14258_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__clkbuf_1
X_19233_ _05693_ _05970_ _05971_ _05696_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a22o_1
X_16445_ registers\[16\]\[10\] registers\[17\]\[10\] registers\[18\]\[10\] registers\[19\]\[10\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14949_ sky130_fd_sc_hd__mux4_1
XFILLER_189_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32491_ clknet_leaf_421_CLK _00605_ VGND VGND VPWR VPWR registers\[60\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_76_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34230_ clknet_leaf_342_CLK _02344_ VGND VGND VPWR VPWR registers\[33\]\[40\] sky130_fd_sc_hd__dfxtp_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19164_ _05688_ _05903_ _05904_ _05691_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__a22o_1
X_31442_ _14222_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__clkbuf_1
X_16376_ registers\[28\]\[8\] registers\[29\]\[8\] registers\[30\]\[8\] registers\[31\]\[8\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14882_ sky130_fd_sc_hd__mux4_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18115_ _04880_ _04883_ _04630_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__o21ba_1
XFILLER_9_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34161_ clknet_leaf_355_CLK _02275_ VGND VGND VPWR VPWR registers\[34\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_31373_ registers\[7\]\[46\] net41 _14179_ VGND VGND VPWR VPWR _14186_ sky130_fd_sc_hd__mux2_1
X_19095_ _05833_ _05836_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__o21ba_1
X_33112_ clknet_leaf_51_CLK _01226_ VGND VGND VPWR VPWR registers\[50\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_30324_ _13633_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__clkbuf_1
X_18046_ registers\[52\]\[56\] registers\[53\]\[56\] registers\[54\]\[56\] registers\[55\]\[56\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__mux4_1
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34092_ clknet_leaf_322_CLK _02206_ VGND VGND VPWR VPWR registers\[35\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33043_ clknet_leaf_74_CLK _01157_ VGND VGND VPWR VPWR registers\[51\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30255_ _13597_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30186_ registers\[16\]\[60\] _13060_ _13494_ VGND VGND VPWR VPWR _13561_ sky130_fd_sc_hd__mux2_1
X_19997_ registers\[52\]\[46\] registers\[53\]\[46\] registers\[54\]\[46\] registers\[55\]\[46\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__mux4_1
XFILLER_99_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18948_ registers\[4\]\[16\] registers\[5\]\[16\] registers\[6\]\[16\] registers\[7\]\[16\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__mux4_1
XANTENNA_1460 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34994_ clknet_leaf_384_CLK _03108_ VGND VGND VPWR VPWR registers\[21\]\[36\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1471 _05328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1482 _06539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1493 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33945_ clknet_leaf_29_CLK _02059_ VGND VGND VPWR VPWR registers\[37\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18879_ registers\[4\]\[14\] registers\[5\]\[14\] registers\[6\]\[14\] registers\[7\]\[14\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__mux4_1
XFILLER_95_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20910_ registers\[40\]\[7\] registers\[41\]\[7\] registers\[42\]\[7\] registers\[43\]\[7\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__mux4_1
XFILLER_228_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33876_ clknet_leaf_120_CLK _01990_ VGND VGND VPWR VPWR registers\[38\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21890_ registers\[24\]\[34\] registers\[25\]\[34\] registers\[26\]\[34\] registers\[27\]\[34\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__mux4_1
XFILLER_81_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20841_ registers\[32\]\[5\] registers\[33\]\[5\] registers\[34\]\[5\] registers\[35\]\[5\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__mux4_1
X_32827_ clknet_leaf_287_CLK _00941_ VGND VGND VPWR VPWR registers\[55\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_35615_ clknet_leaf_485_CLK _03729_ VGND VGND VPWR VPWR registers\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23560_ _09939_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20772_ _07445_ _07452_ _07459_ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__or4_4
X_35546_ clknet_leaf_13_CLK _03660_ VGND VGND VPWR VPWR registers\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_32758_ clknet_leaf_334_CLK _00872_ VGND VGND VPWR VPWR registers\[56\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22511_ _07301_ VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__buf_4
XFILLER_168_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31709_ registers\[59\]\[13\] net5 _14359_ VGND VGND VPWR VPWR _14363_ sky130_fd_sc_hd__mux2_1
X_35477_ clknet_leaf_78_CLK _03591_ VGND VGND VPWR VPWR registers\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23491_ _09577_ registers\[19\]\[30\] _09903_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_67_CLK sky130_fd_sc_hd__clkbuf_16
X_32689_ clknet_leaf_366_CLK _00803_ VGND VGND VPWR VPWR registers\[57\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22442_ _07338_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__clkbuf_4
X_34428_ clknet_leaf_187_CLK _02542_ VGND VGND VPWR VPWR registers\[30\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25230_ _10770_ registers\[51\]\[19\] _10876_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__mux2_1
XFILLER_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25161_ _10845_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22373_ _07300_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__clkbuf_4
X_34359_ clknet_leaf_426_CLK _02473_ VGND VGND VPWR VPWR registers\[31\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24112_ _10234_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21324_ _07929_ _08001_ _08004_ _07932_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__a22o_1
XFILLER_50_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25092_ _10798_ registers\[52\]\[32\] _10794_ VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__mux2_1
XFILLER_164_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28920_ _12864_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24043_ _10197_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36029_ clknet_leaf_288_CLK _04143_ VGND VGND VPWR VPWR registers\[63\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_21255_ registers\[16\]\[16\] registers\[17\]\[16\] registers\[18\]\[16\] registers\[19\]\[16\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__mux4_1
XFILLER_102_1292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20206_ _05049_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__clkbuf_8
XFILLER_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28851_ _11801_ registers\[25\]\[34\] _12823_ VGND VGND VPWR VPWR _12828_ sky130_fd_sc_hd__mux2_1
X_21186_ _07732_ _07869_ _07870_ _07735_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__a22o_1
XFILLER_85_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27802_ registers\[33\]\[49\] _10407_ _12266_ VGND VGND VPWR VPWR _12276_ sky130_fd_sc_hd__mux2_1
X_20137_ registers\[48\]\[50\] registers\[49\]\[50\] registers\[50\]\[50\] registers\[51\]\[50\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux4_1
X_28782_ _11732_ registers\[25\]\[1\] _12790_ VGND VGND VPWR VPWR _12792_ sky130_fd_sc_hd__mux2_1
X_25994_ _11292_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27733_ registers\[33\]\[16\] _10338_ _12233_ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__mux2_1
X_20068_ _06776_ _06778_ _06781_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__a22o_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24945_ _10705_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27664_ _12203_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__clkbuf_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24876_ _10657_ VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__clkbuf_8
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29403_ _13149_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_302 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_313 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26615_ _10793_ registers\[41\]\[30\] _11619_ VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__mux2_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _10082_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_324 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27595_ _12167_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_335 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29334_ _13068_ VGND VGND VPWR VPWR _13113_ sky130_fd_sc_hd__buf_4
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26546_ _11582_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_368 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23758_ _10046_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_379 _00093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22709_ registers\[8\]\[58\] registers\[9\]\[58\] registers\[10\]\[58\] registers\[11\]\[58\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__mux4_1
X_29265_ _09672_ registers\[22\]\[7\] _13069_ VGND VGND VPWR VPWR _13077_ sky130_fd_sc_hd__mux2_1
XFILLER_144_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26477_ _11546_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23689_ _10008_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_58_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_58_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28216_ _11841_ registers\[30\]\[53\] _12490_ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__mux2_1
X_16230_ _14564_ VGND VGND VPWR VPWR _14740_ sky130_fd_sc_hd__buf_4
X_25428_ _10990_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29196_ _13032_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16161_ _14570_ _14671_ _14672_ _14582_ VGND VGND VPWR VPWR _14673_ sky130_fd_sc_hd__a22o_1
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28147_ _11771_ registers\[30\]\[20\] _12457_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__mux2_1
X_25359_ _10954_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28078_ _12421_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__clkbuf_1
X_16092_ _14530_ VGND VGND VPWR VPWR _14606_ sky130_fd_sc_hd__buf_4
XFILLER_6_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27029_ _11736_ registers\[38\]\[3\] _11865_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__mux2_1
XFILLER_170_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19920_ _06569_ _06637_ _06638_ _06574_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__a22o_1
XFILLER_155_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30040_ _13484_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__clkbuf_1
X_19851_ registers\[40\]\[42\] registers\[41\]\[42\] registers\[42\]\[42\] registers\[43\]\[42\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__mux4_1
XFILLER_190_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18802_ registers\[56\]\[12\] registers\[57\]\[12\] registers\[58\]\[12\] registers\[59\]\[12\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__mux4_1
XFILLER_123_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19782_ _06498_ _06503_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__o21ba_1
XFILLER_150_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16994_ _14490_ VGND VGND VPWR VPWR _15482_ sky130_fd_sc_hd__buf_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18733_ registers\[8\]\[10\] registers\[9\]\[10\] registers\[10\]\[10\] registers\[11\]\[10\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__mux4_1
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31991_ clknet_leaf_23_CLK _00163_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_1
XTAP_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33730_ clknet_leaf_249_CLK _01844_ VGND VGND VPWR VPWR registers\[41\]\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18664_ registers\[8\]\[8\] registers\[9\]\[8\] registers\[10\]\[8\] registers\[11\]\[8\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__mux4_1
X_30942_ _13959_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _04395_ _04398_ _04301_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__o21ba_1
X_33661_ clknet_leaf_274_CLK _01775_ VGND VGND VPWR VPWR registers\[42\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_30873_ _13923_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__clkbuf_1
X_18595_ registers\[4\]\[6\] registers\[5\]\[6\] registers\[6\]\[6\] registers\[7\]\[6\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__mux4_1
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35400_ clknet_leaf_156_CLK _03514_ VGND VGND VPWR VPWR registers\[15\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32612_ clknet_leaf_441_CLK _00726_ VGND VGND VPWR VPWR registers\[58\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17546_ _04310_ _04317_ _04324_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or4_1
X_33592_ clknet_leaf_340_CLK _01706_ VGND VGND VPWR VPWR registers\[43\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35331_ clknet_leaf_223_CLK _03445_ VGND VGND VPWR VPWR registers\[16\]\[53\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_880 _09538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_891 _09634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32543_ clknet_leaf_470_CLK _00657_ VGND VGND VPWR VPWR registers\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_17477_ _14548_ VGND VGND VPWR VPWR _15951_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_49_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19216_ registers\[36\]\[24\] registers\[37\]\[24\] registers\[38\]\[24\] registers\[39\]\[24\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__mux4_1
Xclkbuf_6_53__f_CLK clknet_5_26_0_CLK VGND VGND VPWR VPWR clknet_6_53__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_35262_ clknet_leaf_190_CLK _03376_ VGND VGND VPWR VPWR registers\[17\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_16428_ registers\[52\]\[10\] registers\[53\]\[10\] registers\[54\]\[10\] registers\[55\]\[10\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14932_ sky130_fd_sc_hd__mux4_1
X_32474_ clknet_leaf_66_CLK _00588_ VGND VGND VPWR VPWR registers\[60\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34213_ clknet_leaf_56_CLK _02327_ VGND VGND VPWR VPWR registers\[33\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_31425_ _14213_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19147_ _05049_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__clkbuf_4
X_16359_ registers\[60\]\[8\] registers\[61\]\[8\] registers\[62\]\[8\] registers\[63\]\[8\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _14865_ sky130_fd_sc_hd__mux4_1
X_35193_ clknet_leaf_310_CLK _03307_ VGND VGND VPWR VPWR registers\[18\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34144_ clknet_leaf_25_CLK _02258_ VGND VGND VPWR VPWR registers\[34\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31356_ registers\[7\]\[38\] net32 _14168_ VGND VGND VPWR VPWR _14177_ sky130_fd_sc_hd__mux2_1
X_19078_ registers\[48\]\[20\] registers\[49\]\[20\] registers\[50\]\[20\] registers\[51\]\[20\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__mux4_1
X_30307_ registers\[15\]\[53\] _13046_ _13621_ VGND VGND VPWR VPWR _13625_ sky130_fd_sc_hd__mux2_1
X_18029_ registers\[28\]\[55\] registers\[29\]\[55\] registers\[30\]\[55\] registers\[31\]\[55\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__mux4_1
XFILLER_173_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34075_ clknet_leaf_18_CLK _02189_ VGND VGND VPWR VPWR registers\[35\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31287_ registers\[7\]\[5\] net56 _14135_ VGND VGND VPWR VPWR _14141_ sky130_fd_sc_hd__mux2_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33026_ clknet_leaf_263_CLK _01140_ VGND VGND VPWR VPWR registers\[52\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_21040_ _07586_ _07727_ _07728_ _07589_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__a22o_1
XFILLER_125_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30238_ registers\[15\]\[20\] _12976_ _13588_ VGND VGND VPWR VPWR _13589_ sky130_fd_sc_hd__mux2_1
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30169_ _13552_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34977_ clknet_leaf_489_CLK _03091_ VGND VGND VPWR VPWR registers\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_22991_ net30 VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1290 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24730_ _10592_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
X_33928_ clknet_leaf_237_CLK _02042_ VGND VGND VPWR VPWR registers\[38\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_21942_ _07331_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__clkbuf_8
XFILLER_243_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21873_ registers\[56\]\[34\] registers\[57\]\[34\] registers\[58\]\[34\] registers\[59\]\[34\]
+ _08537_ _08327_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__mux4_1
X_24661_ _09592_ registers\[55\]\[37\] _10547_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__mux2_1
X_33859_ clknet_leaf_225_CLK _01973_ VGND VGND VPWR VPWR registers\[3\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26400_ _10850_ registers\[43\]\[57\] _11498_ VGND VGND VPWR VPWR _11506_ sky130_fd_sc_hd__mux2_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20824_ _07343_ _07517_ _07518_ _07353_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__a22o_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23612_ _09968_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27380_ _12053_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__clkbuf_1
X_24592_ _09523_ registers\[55\]\[4\] _10514_ VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__mux2_1
XFILLER_35_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26331_ _10781_ registers\[43\]\[24\] _11465_ VGND VGND VPWR VPWR _11470_ sky130_fd_sc_hd__mux2_1
X_23543_ _09630_ registers\[19\]\[55\] _09925_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__mux2_1
X_35529_ clknet_leaf_160_CLK _03643_ VGND VGND VPWR VPWR registers\[13\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20755_ _07448_ _07451_ _07339_ _07341_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__o211a_1
XFILLER_145_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29050_ _12932_ VGND VGND VPWR VPWR _12933_ sky130_fd_sc_hd__buf_8
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26262_ _11433_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
X_23474_ _09561_ registers\[19\]\[22\] _09892_ VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__mux2_1
X_20686_ _07294_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__buf_12
XFILLER_126_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28001_ _11761_ registers\[31\]\[15\] _12375_ VGND VGND VPWR VPWR _12381_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22425_ _09074_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25213_ _10877_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26193_ _11397_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22356_ _08805_ _09005_ _09006_ _08810_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__a22o_1
X_25144_ _10833_ registers\[52\]\[49\] _10815_ VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__mux2_1
XFILLER_137_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21307_ registers\[48\]\[18\] registers\[49\]\[18\] registers\[50\]\[18\] registers\[51\]\[18\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__mux4_1
XFILLER_178_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29952_ _13438_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__clkbuf_1
X_25075_ net20 VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__buf_2
X_22287_ registers\[44\]\[46\] registers\[45\]\[46\] registers\[46\]\[46\] registers\[47\]\[46\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__mux4_1
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28903_ _11853_ registers\[25\]\[59\] _12845_ VGND VGND VPWR VPWR _12855_ sky130_fd_sc_hd__mux2_1
X_24026_ _10188_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21238_ registers\[52\]\[16\] registers\[53\]\[16\] registers\[54\]\[16\] registers\[55\]\[16\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__mux4_1
X_29883_ registers\[18\]\[44\] _13027_ _13397_ VGND VGND VPWR VPWR _13402_ sky130_fd_sc_hd__mux2_1
XFILLER_215_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28834_ _11784_ registers\[25\]\[26\] _12812_ VGND VGND VPWR VPWR _12819_ sky130_fd_sc_hd__mux2_1
XFILLER_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21169_ _07640_ _07852_ _07853_ _07646_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__a22o_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28765_ _12782_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25977_ _11283_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27716_ registers\[33\]\[8\] _10321_ _12222_ VGND VGND VPWR VPWR _12231_ sky130_fd_sc_hd__mux2_1
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24928_ _10696_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28696_ _12746_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__clkbuf_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27647_ _12194_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__clkbuf_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_110 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24859_ _10660_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_121 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17400_ _15876_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_143 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _05080_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__buf_12
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27578_ _12158_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_154 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29317_ _13104_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_187 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17331_ registers\[40\]\[36\] registers\[41\]\[36\] registers\[42\]\[36\] registers\[43\]\[36\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15809_ sky130_fd_sc_hd__mux4_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26529_ _10844_ registers\[42\]\[54\] _11569_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__mux2_1
XANTENNA_198 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29248_ _13067_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17262_ _15739_ _15742_ _15645_ VGND VGND VPWR VPWR _15743_ sky130_fd_sc_hd__o21ba_1
XFILLER_35_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19001_ _05742_ _05745_ _05475_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__o21ba_1
XFILLER_179_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16213_ _14529_ VGND VGND VPWR VPWR _14723_ sky130_fd_sc_hd__buf_6
XFILLER_128_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17193_ _15654_ _15661_ _15668_ _15675_ VGND VGND VPWR VPWR _15676_ sky130_fd_sc_hd__or4_4
X_29179_ net36 VGND VGND VPWR VPWR _13021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31210_ _14100_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__clkbuf_1
X_16144_ registers\[44\]\[2\] registers\[45\]\[2\] registers\[46\]\[2\] registers\[47\]\[2\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14656_ sky130_fd_sc_hd__mux4_1
XFILLER_154_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32190_ clknet_leaf_462_CLK _00304_ VGND VGND VPWR VPWR registers\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31141_ _14063_ VGND VGND VPWR VPWR _14064_ sky130_fd_sc_hd__buf_4
X_16075_ _14576_ VGND VGND VPWR VPWR _14589_ sky130_fd_sc_hd__buf_6
XFILLER_143_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19903_ _05067_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__buf_6
X_31072_ registers\[0\]\[31\] _13000_ _14026_ VGND VGND VPWR VPWR _14028_ sky130_fd_sc_hd__mux2_1
XFILLER_216_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30023_ _13475_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__clkbuf_1
X_34900_ clknet_leaf_98_CLK _03014_ VGND VGND VPWR VPWR registers\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19834_ _06374_ _06554_ _06555_ _06377_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__a22o_1
XFILLER_190_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35880_ clknet_leaf_401_CLK _03994_ VGND VGND VPWR VPWR registers\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34831_ clknet_leaf_116_CLK _02945_ VGND VGND VPWR VPWR registers\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16977_ _15465_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
X_19765_ registers\[16\]\[39\] registers\[17\]\[39\] registers\[18\]\[39\] registers\[19\]\[39\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__mux4_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 DW[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_8
XFILLER_42_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18716_ _05197_ _05467_ _05468_ _05202_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__a22o_1
X_34762_ clknet_leaf_152_CLK _02876_ VGND VGND VPWR VPWR registers\[25\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_702 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ registers\[20\]\[37\] registers\[21\]\[37\] registers\[22\]\[37\] registers\[23\]\[37\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__mux4_1
X_31974_ clknet_leaf_6_CLK _00144_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18647_ _05204_ _05400_ _05401_ _05207_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__a22o_1
X_30925_ _13950_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__clkbuf_1
X_33713_ clknet_leaf_361_CLK _01827_ VGND VGND VPWR VPWR registers\[41\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_34693_ clknet_leaf_220_CLK _02807_ VGND VGND VPWR VPWR registers\[26\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30856_ _09813_ registers\[11\]\[57\] _13906_ VGND VGND VPWR VPWR _13914_ sky130_fd_sc_hd__mux2_1
X_18578_ _05331_ _05334_ _05074_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__o21ba_2
XFILLER_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33644_ clknet_leaf_330_CLK _01758_ VGND VGND VPWR VPWR registers\[42\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17529_ registers\[52\]\[41\] registers\[53\]\[41\] registers\[54\]\[41\] registers\[55\]\[41\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__mux4_1
X_33575_ clknet_leaf_430_CLK _01689_ VGND VGND VPWR VPWR registers\[43\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30787_ _09740_ registers\[11\]\[24\] _13873_ VGND VGND VPWR VPWR _13878_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20540_ registers\[20\]\[62\] registers\[21\]\[62\] registers\[22\]\[62\] registers\[23\]\[62\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__mux4_1
X_32526_ clknet_leaf_139_CLK _00640_ VGND VGND VPWR VPWR registers\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35314_ clknet_leaf_416_CLK _03428_ VGND VGND VPWR VPWR registers\[16\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20471_ _05040_ _07172_ _07173_ _05050_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__a22o_1
X_32457_ clknet_leaf_214_CLK _00571_ VGND VGND VPWR VPWR registers\[29\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_35245_ clknet_leaf_397_CLK _03359_ VGND VGND VPWR VPWR registers\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_22210_ registers\[16\]\[43\] registers\[17\]\[43\] registers\[18\]\[43\] registers\[19\]\[43\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__mux4_1
X_31408_ registers\[7\]\[63\] net60 _14134_ VGND VGND VPWR VPWR _14204_ sky130_fd_sc_hd__mux2_1
X_35176_ clknet_leaf_405_CLK _03290_ VGND VGND VPWR VPWR registers\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_23190_ _09725_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32388_ clknet_leaf_202_CLK _00502_ VGND VGND VPWR VPWR registers\[61\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34127_ clknet_leaf_131_CLK _02241_ VGND VGND VPWR VPWR registers\[34\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22141_ _08761_ _08797_ _08798_ _08764_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__a22o_1
X_31339_ _14134_ VGND VGND VPWR VPWR _14168_ sky130_fd_sc_hd__buf_6
XFILLER_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34058_ clknet_leaf_159_CLK _02172_ VGND VGND VPWR VPWR registers\[36\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_22072_ _08731_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__buf_6
XFILLER_82_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21023_ _07705_ _07710_ _07711_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__o21ba_1
X_25900_ _11243_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
X_33009_ clknet_leaf_367_CLK _01123_ VGND VGND VPWR VPWR registers\[52\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26880_ _11768_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25831_ _10821_ registers\[47\]\[43\] _11203_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__mux2_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28550_ _12669_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__clkbuf_1
X_25762_ _10751_ registers\[47\]\[10\] _11170_ VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__mux2_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22974_ _09577_ registers\[62\]\[30\] _09578_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__mux2_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27501_ _11803_ registers\[35\]\[35\] _12111_ VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__mux2_1
X_24713_ _09644_ registers\[55\]\[62\] _10513_ VGND VGND VPWR VPWR _10582_ sky130_fd_sc_hd__mux2_1
XFILLER_16_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28481_ _12633_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__clkbuf_1
X_21925_ registers\[28\]\[35\] registers\[29\]\[35\] registers\[30\]\[35\] registers\[31\]\[35\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__mux4_1
XFILLER_216_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25693_ _11133_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_924 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27432_ _11734_ registers\[35\]\[2\] _12078_ VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__mux2_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24644_ _09575_ registers\[55\]\[29\] _10536_ VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__mux2_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21856_ registers\[24\]\[33\] registers\[25\]\[33\] registers\[26\]\[33\] registers\[27\]\[33\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__mux4_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20807_ registers\[32\]\[4\] registers\[33\]\[4\] registers\[34\]\[4\] registers\[35\]\[4\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__mux4_1
XFILLER_180_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27363_ _12044_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__clkbuf_1
X_24575_ _09644_ registers\[56\]\[62\] _10439_ VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__mux2_1
X_21787_ registers\[16\]\[31\] registers\[17\]\[31\] registers\[18\]\[31\] registers\[19\]\[31\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__mux4_1
XFILLER_230_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29102_ registers\[23\]\[16\] _12968_ _12956_ VGND VGND VPWR VPWR _12969_ sky130_fd_sc_hd__mux2_1
X_26314_ _10764_ registers\[43\]\[16\] _11454_ VGND VGND VPWR VPWR _11461_ sky130_fd_sc_hd__mux2_1
XFILLER_208_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23526_ _09613_ registers\[19\]\[47\] _09914_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__mux2_1
X_27294_ _12008_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20738_ _07281_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__buf_6
XFILLER_141_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29033_ _12923_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26245_ _11424_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20669_ _07355_ _07360_ _07365_ _07367_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__a22o_1
X_23457_ _09544_ registers\[19\]\[14\] _09881_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__mux2_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22408_ _09020_ _09056_ _09057_ _09024_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__a22o_1
XFILLER_136_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26176_ _11388_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23388_ registers\[39\]\[47\] _09791_ _09840_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__mux2_1
X_25127_ _10822_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__clkbuf_1
X_22339_ registers\[0\]\[47\] registers\[1\]\[47\] registers\[2\]\[47\] registers\[3\]\[47\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__mux4_1
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29935_ _13429_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__clkbuf_1
X_25058_ _10775_ registers\[52\]\[21\] _10773_ VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__mux2_1
X_16900_ registers\[4\]\[23\] registers\[5\]\[23\] registers\[6\]\[23\] registers\[7\]\[23\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15391_ sky130_fd_sc_hd__mux4_1
XFILLER_111_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24009_ _10179_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
X_17880_ _04540_ _04654_ _04655_ _04546_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__a22o_1
X_29866_ registers\[18\]\[36\] _13010_ _13386_ VGND VGND VPWR VPWR _13393_ sky130_fd_sc_hd__mux2_1
X_16831_ _15144_ _15322_ _15323_ _15147_ VGND VGND VPWR VPWR _15324_ sky130_fd_sc_hd__a22o_1
X_28817_ _11767_ registers\[25\]\[18\] _12801_ VGND VGND VPWR VPWR _12810_ sky130_fd_sc_hd__mux2_1
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29797_ registers\[18\]\[3\] _12941_ _13353_ VGND VGND VPWR VPWR _13357_ sky130_fd_sc_hd__mux2_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19550_ _05067_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__buf_6
XFILLER_232_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28748_ _12773_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__clkbuf_1
X_16762_ registers\[20\]\[19\] registers\[21\]\[19\] registers\[22\]\[19\] registers\[23\]\[19\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15257_ sky130_fd_sc_hd__mux4_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18501_ registers\[20\]\[3\] registers\[21\]\[3\] registers\[22\]\[3\] registers\[23\]\[3\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__mux4_1
XFILLER_47_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19481_ _06031_ _06211_ _06212_ _06034_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__a22o_1
X_28679_ _12737_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__clkbuf_1
X_16693_ _15168_ _15175_ _15182_ _15189_ VGND VGND VPWR VPWR _15190_ sky130_fd_sc_hd__or4_1
XFILLER_94_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30710_ _13837_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__clkbuf_1
X_18432_ _05150_ _05192_ _05193_ _05160_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31690_ registers\[59\]\[4\] net45 _14348_ VGND VGND VPWR VPWR _14353_ sky130_fd_sc_hd__mux2_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18363_ _05125_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__buf_6
X_30641_ registers\[12\]\[19\] _12974_ _13791_ VGND VGND VPWR VPWR _13801_ sky130_fd_sc_hd__mux2_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17314_ _14504_ VGND VGND VPWR VPWR _15793_ sky130_fd_sc_hd__buf_4
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33360_ clknet_leaf_129_CLK _01474_ VGND VGND VPWR VPWR registers\[46\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30572_ _09797_ registers\[13\]\[50\] _13764_ VGND VGND VPWR VPWR _13765_ sky130_fd_sc_hd__mux2_1
X_18294_ net79 net80 VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__and2_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32311_ clknet_leaf_312_CLK _00425_ VGND VGND VPWR VPWR registers\[19\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_17245_ _15549_ _15724_ _15725_ _15553_ VGND VGND VPWR VPWR _15726_ sky130_fd_sc_hd__a22o_1
X_33291_ clknet_leaf_165_CLK _01405_ VGND VGND VPWR VPWR registers\[48\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35030_ clknet_leaf_97_CLK _03144_ VGND VGND VPWR VPWR registers\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_32242_ clknet_leaf_357_CLK _00356_ VGND VGND VPWR VPWR registers\[39\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17176_ registers\[52\]\[31\] registers\[53\]\[31\] registers\[54\]\[31\] registers\[55\]\[31\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15659_ sky130_fd_sc_hd__mux4_1
XFILLER_143_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16127_ registers\[24\]\[1\] registers\[25\]\[1\] registers\[26\]\[1\] registers\[27\]\[1\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _14640_ sky130_fd_sc_hd__mux4_1
XFILLER_157_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32173_ clknet_leaf_86_CLK _00287_ VGND VGND VPWR VPWR registers\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31124_ registers\[0\]\[56\] _13052_ _14048_ VGND VGND VPWR VPWR _14055_ sky130_fd_sc_hd__mux2_1
X_16058_ _14571_ VGND VGND VPWR VPWR _14572_ sky130_fd_sc_hd__buf_8
XFILLER_192_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31055_ registers\[0\]\[23\] _12983_ _14015_ VGND VGND VPWR VPWR _14019_ sky130_fd_sc_hd__mux2_1
X_35932_ clknet_leaf_478_CLK _04046_ VGND VGND VPWR VPWR registers\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_30006_ _13466_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19817_ _06539_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_2
XFILLER_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35863_ clknet_leaf_82_CLK _03977_ VGND VGND VPWR VPWR registers\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34814_ clknet_leaf_298_CLK _02928_ VGND VGND VPWR VPWR registers\[24\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19748_ _06233_ _06470_ _06471_ _06236_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__a22o_1
X_35794_ clknet_leaf_107_CLK _03908_ VGND VGND VPWR VPWR registers\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34745_ clknet_leaf_310_CLK _02859_ VGND VGND VPWR VPWR registers\[25\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31957_ clknet_leaf_0_CLK _00189_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19679_ registers\[48\]\[37\] registers\[49\]\[37\] registers\[50\]\[37\] registers\[51\]\[37\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__mux4_1
XFILLER_225_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_280_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_280_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21710_ _08376_ _08379_ _08073_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__o21ba_1
X_22690_ registers\[20\]\[57\] registers\[21\]\[57\] registers\[22\]\[57\] registers\[23\]\[57\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__mux4_1
X_30908_ _13941_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31888_ _09762_ registers\[49\]\[34\] _14452_ VGND VGND VPWR VPWR _14457_ sky130_fd_sc_hd__mux2_1
X_34676_ clknet_leaf_413_CLK _02790_ VGND VGND VPWR VPWR registers\[26\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21641_ _08075_ _08311_ _08312_ _08078_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__a22o_1
X_30839_ _09795_ registers\[11\]\[49\] _13895_ VGND VGND VPWR VPWR _13905_ sky130_fd_sc_hd__mux2_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33627_ clknet_leaf_26_CLK _01741_ VGND VGND VPWR VPWR registers\[42\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21572_ registers\[28\]\[25\] registers\[29\]\[25\] registers\[30\]\[25\] registers\[31\]\[25\]
+ _08149_ _08150_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__mux4_1
XFILLER_36_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24360_ net31 VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__buf_4
X_33558_ clknet_leaf_126_CLK _01672_ VGND VGND VPWR VPWR registers\[43\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23311_ registers\[9\]\[52\] _09802_ _09798_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__mux2_1
X_20523_ registers\[48\]\[62\] registers\[49\]\[62\] registers\[50\]\[62\] registers\[51\]\[62\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__mux4_1
XANTENNA_43 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32509_ clknet_leaf_288_CLK _00623_ VGND VGND VPWR VPWR registers\[60\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_24291_ _10335_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
X_33489_ clknet_leaf_130_CLK _01603_ VGND VGND VPWR VPWR registers\[44\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_65 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26030_ _11311_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_87 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20454_ _07157_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__buf_4
XANTENNA_98 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23242_ registers\[9\]\[31\] _09756_ _09754_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__mux2_1
X_35228_ clknet_leaf_5_CLK _03342_ VGND VGND VPWR VPWR registers\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23173_ registers\[9\]\[6\] _09670_ _09709_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__mux2_1
XFILLER_137_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20385_ _07087_ _07090_ _06866_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__o21ba_1
XFILLER_175_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35159_ clknet_leaf_91_CLK _03273_ VGND VGND VPWR VPWR registers\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22124_ _08778_ _08781_ _08740_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__o21ba_1
XTAP_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27981_ _12370_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput150 net150 VGND VGND VPWR VPWR D1[6] sky130_fd_sc_hd__buf_2
XTAP_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput161 net161 VGND VGND VPWR VPWR D2[16] sky130_fd_sc_hd__buf_2
XTAP_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput172 net172 VGND VGND VPWR VPWR D2[26] sky130_fd_sc_hd__buf_2
X_29720_ _13316_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__clkbuf_1
XTAP_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput183 net183 VGND VGND VPWR VPWR D2[36] sky130_fd_sc_hd__buf_2
X_26932_ _11803_ registers\[3\]\[35\] _11793_ VGND VGND VPWR VPWR _11804_ sky130_fd_sc_hd__mux2_1
X_22055_ _08677_ _08713_ _08714_ _08681_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__a22o_1
XTAP_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput194 net194 VGND VGND VPWR VPWR D2[46] sky130_fd_sc_hd__buf_2
XTAP_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ registers\[16\]\[9\] registers\[17\]\[9\] registers\[18\]\[9\] registers\[19\]\[9\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__mux4_1
XFILLER_47_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29651_ _13279_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__clkbuf_1
XTAP_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26863_ net5 VGND VGND VPWR VPWR _11757_ sky130_fd_sc_hd__buf_4
XFILLER_248_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28602_ _11822_ registers\[27\]\[44\] _12692_ VGND VGND VPWR VPWR _12697_ sky130_fd_sc_hd__mux2_1
XFILLER_247_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25814_ _10804_ registers\[47\]\[35\] _11192_ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__mux2_1
X_29582_ _13243_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__clkbuf_1
X_26794_ _11714_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28533_ _11753_ registers\[27\]\[11\] _12659_ VGND VGND VPWR VPWR _12661_ sky130_fd_sc_hd__mux2_1
X_25745_ _10735_ registers\[47\]\[2\] _11159_ VGND VGND VPWR VPWR _11162_ sky130_fd_sc_hd__mux2_1
X_22957_ net18 VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__buf_2
XFILLER_95_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28464_ _12624_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__clkbuf_1
X_21908_ _08326_ _08570_ _08571_ _08332_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__a22o_1
X_25676_ _11124_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22888_ _09520_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27415_ _12071_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24627_ _10537_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21839_ _08501_ _08504_ _08397_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__o21ba_1
X_28395_ _12576_ VGND VGND VPWR VPWR _12588_ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27346_ _12035_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__clkbuf_1
X_24558_ _10499_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23509_ _09596_ registers\[19\]\[39\] _09903_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27277_ _11849_ registers\[37\]\[57\] _11991_ VGND VGND VPWR VPWR _11999_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24489_ _10463_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
X_29016_ _12914_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17030_ _15206_ _15515_ _15516_ _15210_ VGND VGND VPWR VPWR _15517_ sky130_fd_sc_hd__a22o_1
X_26228_ _11415_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26159_ _11379_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18981_ _05688_ _05725_ _05726_ _05691_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__a22o_1
XFILLER_140_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29918_ registers\[18\]\[61\] _13062_ _13352_ VGND VGND VPWR VPWR _13420_ sky130_fd_sc_hd__mux2_1
X_17932_ _14578_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__buf_4
XFILLER_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17863_ _14544_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__buf_4
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29849_ registers\[18\]\[28\] _12993_ _13375_ VGND VGND VPWR VPWR _13384_ sky130_fd_sc_hd__mux2_1
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19602_ registers\[44\]\[35\] registers\[45\]\[35\] registers\[46\]\[35\] registers\[47\]\[35\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__mux4_1
X_16814_ _14991_ _15305_ _15306_ _14996_ VGND VGND VPWR VPWR _15307_ sky130_fd_sc_hd__a22o_1
X_17794_ registers\[40\]\[49\] registers\[41\]\[49\] registers\[42\]\[49\] registers\[43\]\[49\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__mux4_1
X_32860_ clknet_leaf_53_CLK _00974_ VGND VGND VPWR VPWR registers\[54\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31811_ registers\[59\]\[62\] net59 _14347_ VGND VGND VPWR VPWR _14416_ sky130_fd_sc_hd__mux2_1
X_19533_ registers\[40\]\[33\] registers\[41\]\[33\] registers\[42\]\[33\] registers\[43\]\[33\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__mux4_1
X_16745_ registers\[48\]\[19\] registers\[49\]\[19\] registers\[50\]\[19\] registers\[51\]\[19\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15240_ sky130_fd_sc_hd__mux4_1
X_32791_ clknet_leaf_61_CLK _00905_ VGND VGND VPWR VPWR registers\[55\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_262_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_262_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19464_ _06196_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__buf_2
X_34530_ clknet_leaf_473_CLK _02644_ VGND VGND VPWR VPWR registers\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_31742_ registers\[59\]\[29\] net22 _14370_ VGND VGND VPWR VPWR _14380_ sky130_fd_sc_hd__mux2_1
X_16676_ registers\[52\]\[17\] registers\[53\]\[17\] registers\[54\]\[17\] registers\[55\]\[17\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15173_ sky130_fd_sc_hd__mux4_1
XFILLER_222_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18415_ _05077_ _05175_ _05176_ _05086_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a22o_1
XFILLER_61_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31673_ _14343_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34461_ clknet_leaf_10_CLK _02575_ VGND VGND VPWR VPWR registers\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ _05890_ _06127_ _06128_ _05893_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__a22o_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36200_ clknet_leaf_22_CLK _00082_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dfxtp_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33412_ clknet_leaf_251_CLK _01526_ VGND VGND VPWR VPWR registers\[46\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_18346_ _05053_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__buf_6
XFILLER_37_1354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30624_ _13792_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34392_ clknet_leaf_19_CLK _02506_ VGND VGND VPWR VPWR registers\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33343_ clknet_leaf_273_CLK _01457_ VGND VGND VPWR VPWR registers\[47\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_36131_ clknet_leaf_47_CLK _04245_ VGND VGND VPWR VPWR registers\[49\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_18277_ _05039_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30555_ _09780_ registers\[13\]\[42\] _13753_ VGND VGND VPWR VPWR _13756_ sky130_fd_sc_hd__mux2_1
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17228_ registers\[20\]\[32\] registers\[21\]\[32\] registers\[22\]\[32\] registers\[23\]\[32\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15710_ sky130_fd_sc_hd__mux4_1
XFILLER_200_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33274_ clknet_leaf_281_CLK _01388_ VGND VGND VPWR VPWR registers\[48\]\[44\] sky130_fd_sc_hd__dfxtp_1
Xinput30 DW[36] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
X_36062_ clknet_leaf_42_CLK _04176_ VGND VGND VPWR VPWR registers\[59\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30486_ _13719_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__clkbuf_1
Xinput41 DW[46] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_8
Xinput52 DW[56] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_16
XFILLER_200_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput63 DW[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_6
X_32225_ clknet_leaf_215_CLK _00339_ VGND VGND VPWR VPWR registers\[9\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_35013_ clknet_leaf_205_CLK _03127_ VGND VGND VPWR VPWR registers\[21\]\[55\] sky130_fd_sc_hd__dfxtp_1
Xinput74 R2[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17159_ _14610_ VGND VGND VPWR VPWR _15643_ sky130_fd_sc_hd__clkbuf_4
Xinput85 RW[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_6
XFILLER_115_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20170_ _06882_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32156_ clknet_leaf_23_CLK _00270_ VGND VGND VPWR VPWR registers\[39\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31107_ registers\[0\]\[48\] _13035_ _14037_ VGND VGND VPWR VPWR _14046_ sky130_fd_sc_hd__mux2_1
XFILLER_233_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32087_ clknet_leaf_489_CLK _00063_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35915_ clknet_leaf_150_CLK _04029_ VGND VGND VPWR VPWR registers\[7\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_31038_ registers\[0\]\[15\] _12966_ _14004_ VGND VGND VPWR VPWR _14010_ sky130_fd_sc_hd__mux2_1
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35846_ clknet_leaf_216_CLK _03960_ VGND VGND VPWR VPWR registers\[8\]\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23860_ _09535_ registers\[60\]\[10\] _10100_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__mux2_1
XFILLER_111_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_0__f_CLK clknet_5_0_0_CLK VGND VGND VPWR VPWR clknet_6_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_22811_ _07355_ _09447_ _09448_ _07367_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__a22o_1
XFILLER_226_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35777_ clknet_leaf_240_CLK _03891_ VGND VGND VPWR VPWR registers\[0\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_23791_ _09603_ registers\[29\]\[42\] _10061_ VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32989_ clknet_leaf_53_CLK _01103_ VGND VGND VPWR VPWR registers\[52\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_709 _07295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_253_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_253_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25530_ _11046_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__clkbuf_1
X_22742_ registers\[12\]\[59\] registers\[13\]\[59\] registers\[14\]\[59\] registers\[15\]\[59\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__mux4_1
XFILLER_37_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34728_ clknet_leaf_452_CLK _02842_ VGND VGND VPWR VPWR registers\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25461_ _11007_ VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__buf_8
XFILLER_213_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22673_ registers\[48\]\[57\] registers\[49\]\[57\] registers\[50\]\[57\] registers\[51\]\[57\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34659_ clknet_leaf_445_CLK _02773_ VGND VGND VPWR VPWR registers\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27200_ _11771_ registers\[37\]\[20\] _11958_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__mux2_1
XFILLER_240_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24412_ _10417_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28180_ _11805_ registers\[30\]\[36\] _12468_ VGND VGND VPWR VPWR _12475_ sky130_fd_sc_hd__mux2_1
X_21624_ _08290_ _08295_ _08054_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__o21ba_1
X_25392_ _10796_ registers\[50\]\[31\] _10970_ VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__mux2_1
XFILLER_194_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27131_ _11922_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24343_ registers\[57\]\[31\] _10370_ _10368_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21555_ _07983_ _08227_ _08228_ _07989_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__a22o_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20506_ registers\[24\]\[61\] registers\[25\]\[61\] registers\[26\]\[61\] registers\[27\]\[61\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__mux4_1
XFILLER_222_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27062_ _11769_ registers\[38\]\[19\] _11876_ VGND VGND VPWR VPWR _11886_ sky130_fd_sc_hd__mux2_1
X_24274_ registers\[57\]\[9\] _10323_ _10305_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__mux2_1
X_21486_ _08158_ _08161_ _08054_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__o21ba_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26013_ _10733_ registers\[45\]\[1\] _11301_ VGND VGND VPWR VPWR _11303_ sky130_fd_sc_hd__mux2_1
X_20437_ _05149_ _07139_ _07140_ _05159_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__a22o_1
X_23225_ _09745_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23156_ _09704_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__buf_8
X_20368_ registers\[44\]\[57\] registers\[45\]\[57\] registers\[46\]\[57\] registers\[47\]\[57\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__mux4_1
XFILLER_164_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1108 _14559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22107_ _07295_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23087_ _09657_ VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__buf_4
XANTENNA_1119 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27964_ registers\[32\]\[62\] _10434_ _12292_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__mux2_1
XTAP_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ registers\[28\]\[54\] registers\[29\]\[54\] registers\[30\]\[54\] registers\[31\]\[54\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__mux4_1
XTAP_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26915_ net24 VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__buf_4
X_29703_ _13307_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__clkbuf_1
X_22038_ _08695_ _08698_ _08430_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__o21ba_1
XTAP_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27895_ registers\[32\]\[29\] _10365_ _12315_ VGND VGND VPWR VPWR _12325_ sky130_fd_sc_hd__mux2_1
XFILLER_212_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_492_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_492_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_29634_ registers\[20\]\[54\] _13048_ _13266_ VGND VGND VPWR VPWR _13271_ sky130_fd_sc_hd__mux2_1
XTAP_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26846_ _11745_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_1
XTAP_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29565_ registers\[20\]\[21\] _12979_ _13233_ VGND VGND VPWR VPWR _13235_ sky130_fd_sc_hd__mux2_1
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26777_ _11705_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23989_ _09529_ registers\[5\]\[7\] _10161_ VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__mux2_1
XFILLER_44_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_244_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_244_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28516_ _11736_ registers\[27\]\[3\] _12648_ VGND VGND VPWR VPWR _12652_ sky130_fd_sc_hd__mux2_1
X_16530_ registers\[44\]\[13\] registers\[45\]\[13\] registers\[46\]\[13\] registers\[47\]\[13\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15031_ sky130_fd_sc_hd__mux4_1
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25728_ _11151_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29496_ _13198_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16461_ _14648_ _14962_ _14963_ _14653_ VGND VGND VPWR VPWR _14964_ sky130_fd_sc_hd__a22o_1
X_28447_ _12615_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__clkbuf_1
X_25659_ _11115_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18200_ registers\[0\]\[61\] registers\[1\]\[61\] registers\[2\]\[61\] registers\[3\]\[61\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__mux4_1
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19180_ registers\[40\]\[23\] registers\[41\]\[23\] registers\[42\]\[23\] registers\[43\]\[23\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__mux4_1
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28378_ _12579_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__clkbuf_1
X_16392_ registers\[48\]\[9\] registers\[49\]\[9\] registers\[50\]\[9\] registers\[51\]\[9\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _14897_ sky130_fd_sc_hd__mux4_1
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ _04895_ _04898_ _04611_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__o21ba_2
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27329_ _12026_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__clkbuf_1
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18062_ _04829_ _04832_ _04644_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__o21ba_1
X_30340_ _09666_ registers\[14\]\[4\] _13638_ VGND VGND VPWR VPWR _13643_ sky130_fd_sc_hd__mux2_1
XFILLER_184_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17013_ _15497_ _15500_ _15302_ VGND VGND VPWR VPWR _15501_ sky130_fd_sc_hd__o21ba_1
XFILLER_156_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30271_ registers\[15\]\[36\] _13010_ _13599_ VGND VGND VPWR VPWR _13606_ sky130_fd_sc_hd__mux2_1
X_32010_ clknet_leaf_29_CLK _00184_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18964_ registers\[32\]\[17\] registers\[33\]\[17\] registers\[34\]\[17\] registers\[35\]\[17\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__mux4_1
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1620 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1631 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17915_ registers\[48\]\[52\] registers\[49\]\[52\] registers\[50\]\[52\] registers\[51\]\[52\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux4_1
XANTENNA_1642 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1653 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33961_ clknet_leaf_424_CLK _02075_ VGND VGND VPWR VPWR registers\[37\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1664 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18895_ _05540_ _05641_ _05642_ _05545_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__a22o_1
XTAP_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1675 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_483_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_483_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35700_ clknet_leaf_415_CLK _03814_ VGND VGND VPWR VPWR registers\[10\]\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1686 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32912_ clknet_leaf_175_CLK _01026_ VGND VGND VPWR VPWR registers\[53\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17846_ _14571_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_1697 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33892_ clknet_leaf_440_CLK _02006_ VGND VGND VPWR VPWR registers\[38\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35631_ clknet_leaf_376_CLK _03745_ VGND VGND VPWR VPWR registers\[11\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32843_ clknet_leaf_166_CLK _00957_ VGND VGND VPWR VPWR registers\[55\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_17777_ registers\[0\]\[48\] registers\[1\]\[48\] registers\[2\]\[48\] registers\[3\]\[48\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__mux4_1
XFILLER_130_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19516_ registers\[0\]\[32\] registers\[1\]\[32\] registers\[2\]\[32\] registers\[3\]\[32\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux4_1
XFILLER_235_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35562_ clknet_leaf_397_CLK _03676_ VGND VGND VPWR VPWR registers\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_16728_ _14947_ _15222_ _15223_ _14950_ VGND VGND VPWR VPWR _15224_ sky130_fd_sc_hd__a22o_1
X_32774_ clknet_leaf_262_CLK _00888_ VGND VGND VPWR VPWR registers\[56\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34513_ clknet_leaf_101_CLK _02627_ VGND VGND VPWR VPWR registers\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16659_ _14952_ _15155_ _15156_ _14957_ VGND VGND VPWR VPWR _15157_ sky130_fd_sc_hd__a22o_1
X_19447_ _05133_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__clkbuf_4
X_31725_ _14371_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35493_ clknet_leaf_463_CLK _03607_ VGND VGND VPWR VPWR registers\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34444_ clknet_leaf_141_CLK _02558_ VGND VGND VPWR VPWR registers\[30\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_31656_ registers\[63\]\[52\] net48 _14332_ VGND VGND VPWR VPWR _14335_ sky130_fd_sc_hd__mux2_1
XFILLER_179_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19378_ _06107_ _06112_ _05837_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__o21ba_1
XFILLER_37_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30607_ _13783_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__clkbuf_1
X_18329_ _05044_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__buf_12
XFILLER_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34375_ clknet_leaf_206_CLK _02489_ VGND VGND VPWR VPWR registers\[31\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_31587_ _14298_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_1378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36114_ clknet_leaf_74_CLK _04228_ VGND VGND VPWR VPWR registers\[49\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21340_ registers\[44\]\[19\] registers\[45\]\[19\] registers\[46\]\[19\] registers\[47\]\[19\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__mux4_1
X_30538_ _09762_ registers\[13\]\[34\] _13742_ VGND VGND VPWR VPWR _13747_ sky130_fd_sc_hd__mux2_1
X_33326_ clknet_leaf_360_CLK _01440_ VGND VGND VPWR VPWR registers\[47\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36045_ clknet_leaf_169_CLK _04159_ VGND VGND VPWR VPWR registers\[63\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_21271_ _07947_ _07952_ _07711_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__o21ba_1
XFILLER_239_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30469_ _09660_ registers\[13\]\[1\] _13709_ VGND VGND VPWR VPWR _13711_ sky130_fd_sc_hd__mux2_1
X_33257_ clknet_leaf_424_CLK _01371_ VGND VGND VPWR VPWR registers\[48\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20222_ registers\[0\]\[52\] registers\[1\]\[52\] registers\[2\]\[52\] registers\[3\]\[52\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__mux4_1
XFILLER_144_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23010_ net37 VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32208_ clknet_leaf_331_CLK _00322_ VGND VGND VPWR VPWR registers\[9\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_33188_ clknet_leaf_471_CLK _01302_ VGND VGND VPWR VPWR registers\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20153_ _05133_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__buf_2
XFILLER_131_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32139_ clknet_leaf_461_CLK _00057_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24961_ _09619_ registers\[53\]\[50\] _10713_ VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__mux2_1
X_20084_ _06793_ _06798_ _06523_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__o21ba_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26700_ registers\[40\]\[6\] _10317_ _11658_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__mux2_1
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_474_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_474_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _09588_ registers\[60\]\[35\] _10122_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__mux2_1
XFILLER_57_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27680_ registers\[34\]\[55\] _10420_ _12206_ VGND VGND VPWR VPWR _12212_ sky130_fd_sc_hd__mux2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24892_ _10677_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26631_ _10810_ registers\[41\]\[38\] _11619_ VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__mux2_1
XFILLER_79_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23843_ _09519_ registers\[60\]\[2\] _10089_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__mux2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35829_ clknet_leaf_353_CLK _03943_ VGND VGND VPWR VPWR registers\[8\]\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_226_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_226_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_506 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29350_ _13121_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_517 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26562_ _10741_ registers\[41\]\[5\] _11586_ VGND VGND VPWR VPWR _11592_ sky130_fd_sc_hd__mux2_1
XANTENNA_528 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23774_ _09586_ registers\[29\]\[34\] _10050_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__mux2_1
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _07433_ _07672_ _07675_ _07438_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__a22o_1
XANTENNA_539 _00183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28301_ _12538_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__clkbuf_1
X_25513_ _11037_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22725_ registers\[40\]\[59\] registers\[41\]\[59\] registers\[42\]\[59\] registers\[43\]\[59\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__mux4_1
X_29281_ _13085_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26493_ _10808_ registers\[42\]\[37\] _11547_ VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__mux2_1
XFILLER_214_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28232_ _11857_ registers\[30\]\[61\] _12434_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25444_ _10848_ registers\[50\]\[56\] _10992_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__mux2_1
X_22656_ registers\[24\]\[56\] registers\[25\]\[56\] registers\[26\]\[56\] registers\[27\]\[56\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__mux4_1
XFILLER_213_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28163_ _11788_ registers\[30\]\[28\] _12457_ VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__mux2_1
X_21607_ _07379_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__buf_4
XFILLER_55_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25375_ _10779_ registers\[50\]\[23\] _10959_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__mux2_1
XFILLER_90_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22587_ registers\[8\]\[54\] registers\[9\]\[54\] registers\[10\]\[54\] registers\[11\]\[54\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__mux4_1
XFILLER_139_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27114_ _11913_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24326_ net19 VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__buf_4
X_28094_ _12429_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__clkbuf_1
X_21538_ registers\[16\]\[24\] registers\[17\]\[24\] registers\[18\]\[24\] registers\[19\]\[24\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__mux4_1
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27045_ _11877_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__clkbuf_1
X_24257_ _10312_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
X_21469_ registers\[24\]\[22\] registers\[25\]\[22\] registers\[26\]\[22\] registers\[27\]\[22\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__mux4_1
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23208_ _09708_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__buf_4
XFILLER_218_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24188_ _09592_ registers\[58\]\[37\] _10266_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__mux2_1
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23139_ net9 VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__buf_4
XTAP_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28996_ registers\[24\]\[39\] _10386_ _12894_ VGND VGND VPWR VPWR _12904_ sky130_fd_sc_hd__mux2_1
XTAP_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27947_ _12352_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__clkbuf_1
XTAP_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17700_ _14490_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__buf_4
XTAP_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_465_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_465_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _05403_ _05418_ _05427_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or4_4
XFILLER_114_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27878_ _12316_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__clkbuf_1
XTAP_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29617_ registers\[20\]\[46\] _13031_ _13255_ VGND VGND VPWR VPWR _13262_ sky130_fd_sc_hd__mux2_1
X_17631_ registers\[52\]\[44\] registers\[53\]\[44\] registers\[54\]\[44\] registers\[55\]\[44\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__mux4_1
X_26829_ net23 VGND VGND VPWR VPWR _11734_ sky130_fd_sc_hd__clkbuf_4
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_247_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_217_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_217_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17562_ registers\[48\]\[42\] registers\[49\]\[42\] registers\[50\]\[42\] registers\[51\]\[42\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__mux4_1
X_29548_ registers\[20\]\[13\] _12962_ _13222_ VGND VGND VPWR VPWR _13226_ sky130_fd_sc_hd__mux2_1
XFILLER_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19301_ registers\[4\]\[26\] registers\[5\]\[26\] registers\[6\]\[26\] registers\[7\]\[26\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__mux4_1
XFILLER_1_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16513_ registers\[4\]\[12\] registers\[5\]\[12\] registers\[6\]\[12\] registers\[7\]\[12\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15015_ sky130_fd_sc_hd__mux4_1
XFILLER_56_1004 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17493_ _14571_ VGND VGND VPWR VPWR _15967_ sky130_fd_sc_hd__buf_4
XFILLER_210_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29479_ _13189_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31510_ _09791_ registers\[6\]\[47\] _14250_ VGND VGND VPWR VPWR _14258_ sky130_fd_sc_hd__mux2_1
XFILLER_231_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19232_ registers\[4\]\[24\] registers\[5\]\[24\] registers\[6\]\[24\] registers\[7\]\[24\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__mux4_1
XFILLER_32_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16444_ registers\[24\]\[10\] registers\[25\]\[10\] registers\[26\]\[10\] registers\[27\]\[10\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14948_ sky130_fd_sc_hd__mux4_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32490_ clknet_leaf_407_CLK _00604_ VGND VGND VPWR VPWR registers\[60\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19163_ registers\[0\]\[22\] registers\[1\]\[22\] registers\[2\]\[22\] registers\[3\]\[22\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__mux4_1
X_31441_ _09687_ registers\[6\]\[14\] _14217_ VGND VGND VPWR VPWR _14222_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16375_ _14588_ _14879_ _14880_ _14598_ VGND VGND VPWR VPWR _14881_ sky130_fd_sc_hd__a22o_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18114_ _14511_ _04881_ _04882_ _14517_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a22o_1
XFILLER_158_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34160_ clknet_leaf_349_CLK _02274_ VGND VGND VPWR VPWR registers\[34\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_31372_ _14185_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__clkbuf_1
X_19094_ _05133_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__buf_2
XFILLER_160_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30323_ registers\[15\]\[61\] _13062_ _13565_ VGND VGND VPWR VPWR _13633_ sky130_fd_sc_hd__mux2_1
X_18045_ registers\[60\]\[56\] registers\[61\]\[56\] registers\[62\]\[56\] registers\[63\]\[56\]
+ _04755_ _04549_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux4_1
X_33111_ clknet_leaf_68_CLK _01225_ VGND VGND VPWR VPWR registers\[50\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34091_ clknet_leaf_425_CLK _02205_ VGND VGND VPWR VPWR registers\[35\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33042_ clknet_leaf_73_CLK _01156_ VGND VGND VPWR VPWR registers\[51\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_30254_ registers\[15\]\[28\] _12993_ _13588_ VGND VGND VPWR VPWR _13597_ sky130_fd_sc_hd__mux2_1
XFILLER_235_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30185_ _13560_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__clkbuf_1
X_19996_ _05097_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__buf_4
XFILLER_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18947_ registers\[12\]\[16\] registers\[13\]\[16\] registers\[14\]\[16\] registers\[15\]\[16\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__mux4_1
XFILLER_100_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_13__f_CLK clknet_5_6_0_CLK VGND VGND VPWR VPWR clknet_6_13__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_34993_ clknet_leaf_381_CLK _03107_ VGND VGND VPWR VPWR registers\[21\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1450 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1461 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_456_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_456_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_239_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1472 _05328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1483 _06807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33944_ clknet_leaf_31_CLK _02058_ VGND VGND VPWR VPWR registers\[37\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_18878_ registers\[12\]\[14\] registers\[13\]\[14\] registers\[14\]\[14\] registers\[15\]\[14\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__mux4_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1494 _07324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17829_ _14546_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__buf_4
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33875_ clknet_leaf_126_CLK _01989_ VGND VGND VPWR VPWR registers\[38\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_208_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_208_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35614_ clknet_leaf_485_CLK _03728_ VGND VGND VPWR VPWR registers\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_20840_ registers\[40\]\[5\] registers\[41\]\[5\] registers\[42\]\[5\] registers\[43\]\[5\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__mux4_1
X_32826_ clknet_leaf_287_CLK _00940_ VGND VGND VPWR VPWR registers\[55\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35545_ clknet_leaf_13_CLK _03659_ VGND VGND VPWR VPWR registers\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_20771_ _07462_ _07467_ _07399_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__o21ba_1
XFILLER_50_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32757_ clknet_leaf_351_CLK _00871_ VGND VGND VPWR VPWR registers\[56\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22510_ registers\[36\]\[52\] registers\[37\]\[52\] registers\[38\]\[52\] registers\[39\]\[52\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__mux4_1
X_31708_ _14362_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__clkbuf_1
X_35476_ clknet_leaf_81_CLK _03590_ VGND VGND VPWR VPWR registers\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_23490_ _09869_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__buf_4
X_32688_ clknet_leaf_366_CLK _00802_ VGND VGND VPWR VPWR registers\[57\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22441_ _09020_ _09088_ _09089_ _09024_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__a22o_1
X_34427_ clknet_leaf_184_CLK _02541_ VGND VGND VPWR VPWR registers\[30\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31639_ registers\[63\]\[44\] net39 _14321_ VGND VGND VPWR VPWR _14326_ sky130_fd_sc_hd__mux2_1
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25160_ _10844_ registers\[52\]\[54\] _10836_ VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__mux2_1
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22372_ registers\[52\]\[48\] registers\[53\]\[48\] registers\[54\]\[48\] registers\[55\]\[48\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__mux4_1
X_34358_ clknet_leaf_426_CLK _02472_ VGND VGND VPWR VPWR registers\[31\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_24111_ _09510_ registers\[58\]\[0\] _10233_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__mux2_1
X_33309_ clknet_leaf_28_CLK _01423_ VGND VGND VPWR VPWR registers\[47\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_21323_ registers\[4\]\[18\] registers\[5\]\[18\] registers\[6\]\[18\] registers\[7\]\[18\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__mux4_1
XFILLER_11_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25091_ net26 VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__clkbuf_4
X_34289_ clknet_leaf_355_CLK _02403_ VGND VGND VPWR VPWR registers\[32\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_36028_ clknet_leaf_288_CLK _04142_ VGND VGND VPWR VPWR registers\[63\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24042_ _09582_ registers\[5\]\[32\] _10194_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__mux2_1
X_21254_ _07379_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__buf_4
XFILLER_102_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20205_ registers\[32\]\[52\] registers\[33\]\[52\] registers\[34\]\[52\] registers\[35\]\[52\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__mux4_1
X_28850_ _12827_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__clkbuf_1
X_21185_ registers\[16\]\[14\] registers\[17\]\[14\] registers\[18\]\[14\] registers\[19\]\[14\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__mux4_1
XFILLER_143_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20136_ registers\[56\]\[50\] registers\[57\]\[50\] registers\[58\]\[50\] registers\[59\]\[50\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__mux4_1
X_27801_ _12275_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__clkbuf_1
X_28781_ _12791_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25993_ _10848_ registers\[46\]\[56\] _11285_ VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_447_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_447_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27732_ _12239_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__clkbuf_1
X_20067_ _05048_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__clkbuf_4
XFILLER_161_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24944_ _09603_ registers\[53\]\[42\] _10702_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__mux2_1
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27663_ registers\[34\]\[47\] _10403_ _12195_ VGND VGND VPWR VPWR _12203_ sky130_fd_sc_hd__mux2_1
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24875_ _10668_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__clkbuf_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29402_ _09674_ registers\[21\]\[8\] _13140_ VGND VGND VPWR VPWR _13149_ sky130_fd_sc_hd__mux2_1
X_26614_ _11585_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__clkbuf_8
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23826_ _09638_ registers\[29\]\[59\] _10072_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_303 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27594_ registers\[34\]\[14\] _10334_ _12162_ VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__mux2_1
XANTENNA_325 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_336 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_347 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26545_ _10860_ registers\[42\]\[62\] _11513_ VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__mux2_1
X_29333_ _13112_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__clkbuf_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23757_ _09569_ registers\[29\]\[26\] _10039_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__mux2_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _07363_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__buf_4
XANTENNA_369 _00092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22708_ _09345_ _09348_ _09091_ _09092_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__o211a_1
X_29264_ _13076_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26476_ _10791_ registers\[42\]\[29\] _11536_ VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__mux2_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23688_ registers\[61\]\[59\] _09817_ _09998_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__mux2_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28215_ _12493_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25427_ _10831_ registers\[50\]\[48\] _10981_ VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__mux2_1
X_22639_ registers\[36\]\[56\] registers\[37\]\[56\] registers\[38\]\[56\] registers\[39\]\[56\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__mux4_1
X_29195_ registers\[23\]\[46\] _13031_ _13019_ VGND VGND VPWR VPWR _13032_ sky130_fd_sc_hd__mux2_1
XFILLER_142_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16160_ registers\[4\]\[2\] registers\[5\]\[2\] registers\[6\]\[2\] registers\[7\]\[2\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14672_ sky130_fd_sc_hd__mux4_1
X_28146_ _12434_ VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__buf_4
X_25358_ _10762_ registers\[50\]\[15\] _10948_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24309_ registers\[57\]\[20\] _10346_ _10347_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__mux2_1
X_16091_ registers\[28\]\[0\] registers\[29\]\[0\] registers\[30\]\[0\] registers\[31\]\[0\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _14605_ sky130_fd_sc_hd__mux4_1
X_28077_ _11837_ registers\[31\]\[51\] _12419_ VGND VGND VPWR VPWR _12421_ sky130_fd_sc_hd__mux2_1
XFILLER_86_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25289_ _10829_ registers\[51\]\[47\] _10909_ VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__mux2_1
XFILLER_170_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_851 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27028_ _11868_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19850_ _05045_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18801_ _05546_ _05551_ _05475_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__o21ba_1
X_19781_ _05073_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__buf_2
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28979_ _12895_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__clkbuf_1
X_16993_ _15475_ _15480_ _15277_ _15278_ VGND VGND VPWR VPWR _15481_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_438_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_438_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18732_ _05479_ _05482_ _05483_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__o211a_2
XTAP_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31990_ clknet_leaf_23_CLK _00162_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ _05411_ _05417_ _05103_ _05105_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__o211a_1
X_30941_ registers\[10\]\[33\] _13004_ _13955_ VGND VGND VPWR VPWR _13959_ sky130_fd_sc_hd__mux2_1
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _04294_ _04396_ _04397_ _04299_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a22o_1
X_33660_ clknet_leaf_277_CLK _01774_ VGND VGND VPWR VPWR registers\[42\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30872_ registers\[10\]\[0\] _12931_ _13922_ VGND VGND VPWR VPWR _13923_ sky130_fd_sc_hd__mux2_1
X_18594_ registers\[12\]\[6\] registers\[13\]\[6\] registers\[14\]\[6\] registers\[15\]\[6\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__mux4_1
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32611_ clknet_leaf_443_CLK _00725_ VGND VGND VPWR VPWR registers\[58\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17545_ _04327_ _04330_ _04301_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__o21ba_1
XFILLER_17_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33591_ clknet_leaf_341_CLK _01705_ VGND VGND VPWR VPWR registers\[43\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_870 _09480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35330_ clknet_leaf_223_CLK _03444_ VGND VGND VPWR VPWR registers\[16\]\[52\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_881 _09538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_892 _09634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17476_ _14546_ VGND VGND VPWR VPWR _15950_ sky130_fd_sc_hd__buf_4
X_32542_ clknet_leaf_481_CLK _00656_ VGND VGND VPWR VPWR registers\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19215_ registers\[44\]\[24\] registers\[45\]\[24\] registers\[46\]\[24\] registers\[47\]\[24\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__mux4_1
X_35261_ clknet_leaf_190_CLK _03375_ VGND VGND VPWR VPWR registers\[17\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_16427_ registers\[60\]\[10\] registers\[61\]\[10\] registers\[62\]\[10\] registers\[63\]\[10\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _14931_ sky130_fd_sc_hd__mux4_1
X_32473_ clknet_leaf_62_CLK _00587_ VGND VGND VPWR VPWR registers\[60\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34212_ clknet_leaf_56_CLK _02326_ VGND VGND VPWR VPWR registers\[33\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_31424_ _09670_ registers\[6\]\[6\] _14206_ VGND VGND VPWR VPWR _14213_ sky130_fd_sc_hd__mux2_1
X_16358_ _14543_ VGND VGND VPWR VPWR _14864_ sky130_fd_sc_hd__buf_4
XFILLER_34_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19146_ registers\[32\]\[22\] registers\[33\]\[22\] registers\[34\]\[22\] registers\[35\]\[22\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__mux4_1
XFILLER_203_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35192_ clknet_leaf_428_CLK _03306_ VGND VGND VPWR VPWR registers\[18\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31355_ _14176_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__clkbuf_1
X_34143_ clknet_leaf_16_CLK _02257_ VGND VGND VPWR VPWR registers\[34\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_16289_ registers\[8\]\[6\] registers\[9\]\[6\] registers\[10\]\[6\] registers\[11\]\[6\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14797_ sky130_fd_sc_hd__mux4_1
XFILLER_117_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19077_ registers\[56\]\[20\] registers\[57\]\[20\] registers\[58\]\[20\] registers\[59\]\[20\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__mux4_1
XFILLER_117_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30306_ _13624_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__clkbuf_1
X_18028_ _04632_ _04798_ _04799_ _04635_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__a22o_1
XFILLER_246_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31286_ _14140_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34074_ clknet_leaf_18_CLK _02188_ VGND VGND VPWR VPWR registers\[35\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_33025_ clknet_leaf_267_CLK _01139_ VGND VGND VPWR VPWR registers\[52\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_30237_ _13565_ VGND VGND VPWR VPWR _13588_ sky130_fd_sc_hd__buf_4
XFILLER_114_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30168_ registers\[16\]\[51\] _13042_ _13550_ VGND VGND VPWR VPWR _13552_ sky130_fd_sc_hd__mux2_1
XFILLER_140_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19979_ registers\[20\]\[45\] registers\[21\]\[45\] registers\[22\]\[45\] registers\[23\]\[45\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__mux4_1
XFILLER_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_429_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_429_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22990_ _09589_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
X_34976_ clknet_leaf_490_CLK _03090_ VGND VGND VPWR VPWR registers\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_30099_ _13515_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1280 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1291 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33927_ clknet_leaf_236_CLK _02041_ VGND VGND VPWR VPWR registers\[38\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_21941_ registers\[60\]\[36\] registers\[61\]\[36\] registers\[62\]\[36\] registers\[63\]\[36\]
+ _08541_ _08335_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__mux4_1
XFILLER_132_1286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24660_ _10554_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33858_ clknet_leaf_225_CLK _01972_ VGND VGND VPWR VPWR registers\[3\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_21872_ _07314_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__buf_6
XFILLER_167_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ registers\[61\]\[22\] _09717_ _09965_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__mux2_1
X_20823_ registers\[0\]\[4\] registers\[1\]\[4\] registers\[2\]\[4\] registers\[3\]\[4\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__mux4_1
X_32809_ clknet_leaf_423_CLK _00923_ VGND VGND VPWR VPWR registers\[55\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_24591_ _10518_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
X_33789_ clknet_leaf_274_CLK _01903_ VGND VGND VPWR VPWR registers\[40\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26330_ _11469_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
X_23542_ _09930_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
X_35528_ clknet_leaf_155_CLK _03642_ VGND VGND VPWR VPWR registers\[13\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20754_ _07325_ _07449_ _07450_ _07336_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__a22o_1
X_26261_ _10846_ registers\[44\]\[55\] _11427_ VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__mux2_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35459_ clknet_leaf_227_CLK _03573_ VGND VGND VPWR VPWR registers\[14\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23473_ _09894_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20685_ _07373_ _07376_ _07381_ _07383_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__a22o_1
XFILLER_138_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28000_ _12380_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__clkbuf_1
X_25212_ _10751_ registers\[51\]\[10\] _10876_ VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__mux2_1
X_22424_ _09052_ _09059_ _09066_ _09073_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__or4_4
X_26192_ _10777_ registers\[44\]\[22\] _11394_ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__mux2_1
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25143_ net44 VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__buf_2
X_22355_ registers\[32\]\[48\] registers\[33\]\[48\] registers\[34\]\[48\] registers\[35\]\[48\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__mux4_1
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21306_ _07281_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__clkbuf_4
X_29951_ registers\[17\]\[12\] _12960_ _13435_ VGND VGND VPWR VPWR _13438_ sky130_fd_sc_hd__mux2_1
X_25074_ _10786_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
X_22286_ _08805_ _08937_ _08938_ _08810_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__a22o_1
XFILLER_219_1431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28902_ _12854_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__clkbuf_1
X_24025_ _09565_ registers\[5\]\[24\] _10183_ VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__mux2_1
X_21237_ _07333_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__buf_4
X_29882_ _13401_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28833_ _12818_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21168_ registers\[48\]\[14\] registers\[49\]\[14\] registers\[50\]\[14\] registers\[51\]\[14\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20119_ _06525_ _06831_ _06832_ _06528_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__a22o_1
X_28764_ _11849_ registers\[26\]\[57\] _12774_ VGND VGND VPWR VPWR _12782_ sky130_fd_sc_hd__mux2_1
X_25976_ _10831_ registers\[46\]\[48\] _11274_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__mux2_1
X_21099_ _07366_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__clkbuf_4
X_27715_ _12230_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__clkbuf_1
X_24927_ _09586_ registers\[53\]\[34\] _10691_ VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__mux2_1
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28695_ _11780_ registers\[26\]\[24\] _12741_ VGND VGND VPWR VPWR _12746_ sky130_fd_sc_hd__mux2_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24858_ _09517_ registers\[53\]\[1\] _10658_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__mux2_1
XANTENNA_100 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27646_ registers\[34\]\[39\] _10386_ _12184_ VGND VGND VPWR VPWR _12194_ sky130_fd_sc_hd__mux2_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23809_ _10073_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27577_ registers\[34\]\[6\] _10317_ _12151_ VGND VGND VPWR VPWR _12158_ sky130_fd_sc_hd__mux2_1
XANTENNA_144 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24789_ _10623_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_166 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _15808_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__clkbuf_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26528_ _11573_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_177 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29316_ _09756_ registers\[22\]\[31\] _13102_ VGND VGND VPWR VPWR _13104_ sky130_fd_sc_hd__mux2_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_188 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17261_ _15638_ _15740_ _15741_ _15643_ VGND VGND VPWR VPWR _15742_ sky130_fd_sc_hd__a22o_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29247_ registers\[23\]\[63\] _13066_ _12934_ VGND VGND VPWR VPWR _13067_ sky130_fd_sc_hd__mux2_1
XFILLER_198_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26459_ _11537_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16212_ _14718_ _14721_ _14525_ VGND VGND VPWR VPWR _14722_ sky130_fd_sc_hd__o21ba_1
XFILLER_202_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19000_ _05547_ _05743_ _05744_ _05550_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29178_ _13020_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _15671_ _15674_ _15645_ VGND VGND VPWR VPWR _15675_ sky130_fd_sc_hd__o21ba_1
XFILLER_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16143_ _14510_ VGND VGND VPWR VPWR _14655_ sky130_fd_sc_hd__buf_6
X_28129_ _12448_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31140_ _09705_ _11084_ VGND VGND VPWR VPWR _14063_ sky130_fd_sc_hd__nor2_8
X_16074_ _14587_ VGND VGND VPWR VPWR _14588_ sky130_fd_sc_hd__buf_4
XFILLER_6_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19902_ _06374_ _06620_ _06621_ _06377_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__a22o_1
X_31071_ _14027_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30022_ registers\[17\]\[46\] _13031_ _13468_ VGND VGND VPWR VPWR _13475_ sky130_fd_sc_hd__mux2_1
X_19833_ registers\[0\]\[41\] registers\[1\]\[41\] registers\[2\]\[41\] registers\[3\]\[41\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__mux4_1
XFILLER_29_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34830_ clknet_leaf_116_CLK _02944_ VGND VGND VPWR VPWR registers\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19764_ registers\[24\]\[39\] registers\[25\]\[39\] registers\[26\]\[39\] registers\[27\]\[39\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__mux4_1
X_16976_ _15441_ _15448_ _15457_ _15464_ VGND VGND VPWR VPWR _15465_ sky130_fd_sc_hd__or4_4
XFILLER_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18715_ registers\[32\]\[10\] registers\[33\]\[10\] registers\[34\]\[10\] registers\[35\]\[10\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__mux4_1
X_34761_ clknet_leaf_220_CLK _02875_ VGND VGND VPWR VPWR registers\[25\]\[59\] sky130_fd_sc_hd__dfxtp_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 DW[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_8
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31973_ clknet_leaf_6_CLK _00143_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
X_19695_ registers\[28\]\[37\] registers\[29\]\[37\] registers\[30\]\[37\] registers\[31\]\[37\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__mux4_1
XFILLER_225_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33712_ clknet_leaf_347_CLK _01826_ VGND VGND VPWR VPWR registers\[41\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18646_ registers\[36\]\[8\] registers\[37\]\[8\] registers\[38\]\[8\] registers\[39\]\[8\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__mux4_1
X_30924_ registers\[10\]\[25\] _12987_ _13944_ VGND VGND VPWR VPWR _13950_ sky130_fd_sc_hd__mux2_1
X_34692_ clknet_leaf_219_CLK _02806_ VGND VGND VPWR VPWR registers\[26\]\[54\] sky130_fd_sc_hd__dfxtp_1
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33643_ clknet_leaf_428_CLK _01757_ VGND VGND VPWR VPWR registers\[42\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_30855_ _13913_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__clkbuf_1
X_18577_ _05204_ _05332_ _05333_ _05207_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__a22o_1
XFILLER_206_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_196_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17528_ registers\[60\]\[41\] registers\[61\]\[41\] registers\[62\]\[41\] registers\[63\]\[41\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__mux4_1
X_33574_ clknet_leaf_57_CLK _01688_ VGND VGND VPWR VPWR registers\[43\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30786_ _13877_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35313_ clknet_leaf_394_CLK _03427_ VGND VGND VPWR VPWR registers\[16\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_32525_ clknet_leaf_167_CLK _00639_ VGND VGND VPWR VPWR registers\[60\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17459_ _15825_ _15932_ _15933_ _15828_ VGND VGND VPWR VPWR _15934_ sky130_fd_sc_hd__a22o_1
XFILLER_220_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35244_ clknet_leaf_396_CLK _03358_ VGND VGND VPWR VPWR registers\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_20470_ registers\[0\]\[60\] registers\[1\]\[60\] registers\[2\]\[60\] registers\[3\]\[60\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__mux4_1
X_32456_ clknet_leaf_211_CLK _00570_ VGND VGND VPWR VPWR registers\[29\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31407_ _14203_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__clkbuf_1
X_19129_ registers\[12\]\[21\] registers\[13\]\[21\] registers\[14\]\[21\] registers\[15\]\[21\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__mux4_1
X_35175_ clknet_leaf_448_CLK _03289_ VGND VGND VPWR VPWR registers\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_32387_ clknet_leaf_233_CLK _00501_ VGND VGND VPWR VPWR registers\[61\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34126_ clknet_leaf_131_CLK _02240_ VGND VGND VPWR VPWR registers\[34\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_22140_ registers\[16\]\[41\] registers\[17\]\[41\] registers\[18\]\[41\] registers\[19\]\[41\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__mux4_1
X_31338_ _14167_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34057_ clknet_leaf_261_CLK _02171_ VGND VGND VPWR VPWR registers\[36\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_22071_ _08709_ _08716_ _08723_ _08730_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__or4_1
XFILLER_82_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31269_ registers\[8\]\[61\] net58 _14063_ VGND VGND VPWR VPWR _14131_ sky130_fd_sc_hd__mux2_1
XTAP_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21022_ _07309_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__buf_2
X_33008_ clknet_leaf_367_CLK _01122_ VGND VGND VPWR VPWR registers\[52\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25830_ _11206_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25761_ _11158_ VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__buf_4
X_34959_ clknet_leaf_114_CLK _03073_ VGND VGND VPWR VPWR registers\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_22973_ _09514_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__buf_4
XFILLER_74_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24712_ _10581_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
X_27500_ _12116_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__clkbuf_1
X_28480_ _11834_ registers\[28\]\[50\] _12632_ VGND VGND VPWR VPWR _12633_ sky130_fd_sc_hd__mux2_1
X_21924_ _08418_ _08586_ _08587_ _08421_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__a22o_1
X_25692_ registers\[48\]\[42\] _10393_ _11130_ VGND VGND VPWR VPWR _11133_ sky130_fd_sc_hd__mux2_1
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27431_ _12080_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24643_ _10545_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _08515_ _08520_ _08416_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__o21ba_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_215_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ registers\[40\]\[4\] registers\[41\]\[4\] registers\[42\]\[4\] registers\[43\]\[4\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__mux4_1
X_27362_ registers\[36\]\[33\] _10374_ _12040_ VGND VGND VPWR VPWR _12044_ sky130_fd_sc_hd__mux2_1
X_24574_ _10507_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21786_ registers\[24\]\[31\] registers\[25\]\[31\] registers\[26\]\[31\] registers\[27\]\[31\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__mux4_1
XFILLER_145_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29101_ net8 VGND VGND VPWR VPWR _12968_ sky130_fd_sc_hd__clkbuf_4
X_26313_ _11460_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23525_ _09921_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27293_ registers\[36\]\[0\] _10303_ _12007_ VGND VGND VPWR VPWR _12008_ sky130_fd_sc_hd__mux2_1
X_20737_ _07278_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__buf_6
XFILLER_208_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29032_ registers\[24\]\[56\] _10422_ _12916_ VGND VGND VPWR VPWR _12923_ sky130_fd_sc_hd__mux2_1
X_26244_ _10829_ registers\[44\]\[47\] _11416_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__mux2_1
XFILLER_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23456_ _09885_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__clkbuf_1
X_20668_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22407_ registers\[52\]\[49\] registers\[53\]\[49\] registers\[54\]\[49\] registers\[55\]\[49\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__mux4_1
X_26175_ _10760_ registers\[44\]\[14\] _11383_ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__mux2_1
X_23387_ _09847_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
X_20599_ _07289_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_221_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25126_ _10821_ registers\[52\]\[43\] _10815_ VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__mux2_1
X_22338_ registers\[8\]\[47\] registers\[9\]\[47\] registers\[10\]\[47\] registers\[11\]\[47\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__mux4_1
XFILLER_139_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29934_ registers\[17\]\[4\] _12943_ _13424_ VGND VGND VPWR VPWR _13429_ sky130_fd_sc_hd__mux2_1
XFILLER_124_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25057_ net14 VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22269_ registers\[0\]\[45\] registers\[1\]\[45\] registers\[2\]\[45\] registers\[3\]\[45\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__mux4_1
XFILLER_3_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24008_ _09548_ registers\[5\]\[16\] _10172_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__mux2_1
XFILLER_215_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29865_ _13392_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16830_ registers\[4\]\[21\] registers\[5\]\[21\] registers\[6\]\[21\] registers\[7\]\[21\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15323_ sky130_fd_sc_hd__mux4_1
X_28816_ _12809_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29796_ _13356_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28747_ _11832_ registers\[26\]\[49\] _12763_ VGND VGND VPWR VPWR _12773_ sky130_fd_sc_hd__mux2_1
X_16761_ registers\[28\]\[19\] registers\[29\]\[19\] registers\[30\]\[19\] registers\[31\]\[19\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15256_ sky130_fd_sc_hd__mux4_1
X_25959_ _11229_ VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__buf_4
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18500_ registers\[28\]\[3\] registers\[29\]\[3\] registers\[30\]\[3\] registers\[31\]\[3\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__mux4_1
XFILLER_46_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19480_ registers\[0\]\[31\] registers\[1\]\[31\] registers\[2\]\[31\] registers\[3\]\[31\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__mux4_1
X_16692_ _15185_ _15188_ _14959_ VGND VGND VPWR VPWR _15189_ sky130_fd_sc_hd__o21ba_1
XFILLER_234_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28678_ _11763_ registers\[26\]\[16\] _12730_ VGND VGND VPWR VPWR _12737_ sky130_fd_sc_hd__mux2_1
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18431_ registers\[20\]\[1\] registers\[21\]\[1\] registers\[22\]\[1\] registers\[23\]\[1\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__mux4_1
XFILLER_94_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27629_ _12185_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18362_ _05078_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__buf_12
X_30640_ _13800_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17313_ _14502_ VGND VGND VPWR VPWR _15792_ sky130_fd_sc_hd__buf_6
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30571_ _13708_ VGND VGND VPWR VPWR _13764_ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _05040_ _05047_ _05050_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__a22o_1
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32310_ clknet_leaf_312_CLK _00424_ VGND VGND VPWR VPWR registers\[19\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_17244_ registers\[52\]\[33\] registers\[53\]\[33\] registers\[54\]\[33\] registers\[55\]\[33\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15725_ sky130_fd_sc_hd__mux4_1
X_33290_ clknet_leaf_163_CLK _01404_ VGND VGND VPWR VPWR registers\[48\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17175_ registers\[60\]\[31\] registers\[61\]\[31\] registers\[62\]\[31\] registers\[63\]\[31\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15658_ sky130_fd_sc_hd__mux4_1
X_32241_ clknet_leaf_357_CLK _00355_ VGND VGND VPWR VPWR registers\[39\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16126_ _14635_ _14638_ _14585_ VGND VGND VPWR VPWR _14639_ sky130_fd_sc_hd__o21ba_1
X_32172_ clknet_leaf_79_CLK _00286_ VGND VGND VPWR VPWR registers\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31123_ _14054_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__clkbuf_1
X_16057_ _14492_ VGND VGND VPWR VPWR _14571_ sky130_fd_sc_hd__buf_12
XFILLER_170_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31054_ _14018_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__clkbuf_1
X_35931_ clknet_leaf_476_CLK _04045_ VGND VGND VPWR VPWR registers\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30005_ registers\[17\]\[38\] _13014_ _13457_ VGND VGND VPWR VPWR _13466_ sky130_fd_sc_hd__mux2_1
XFILLER_243_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19816_ _06505_ _06514_ _06524_ _06538_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__or4_4
X_35862_ clknet_leaf_69_CLK _03976_ VGND VGND VPWR VPWR registers\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34813_ clknet_leaf_306_CLK _02927_ VGND VGND VPWR VPWR registers\[24\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_19747_ registers\[36\]\[39\] registers\[37\]\[39\] registers\[38\]\[39\] registers\[39\]\[39\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__mux4_1
X_35793_ clknet_leaf_107_CLK _03907_ VGND VGND VPWR VPWR registers\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16959_ _15444_ _15447_ _15277_ _15278_ VGND VGND VPWR VPWR _15448_ sky130_fd_sc_hd__o211a_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34744_ clknet_leaf_426_CLK _02858_ VGND VGND VPWR VPWR registers\[25\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_31956_ clknet_leaf_0_CLK _00188_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_1
X_19678_ registers\[56\]\[37\] registers\[57\]\[37\] registers\[58\]\[37\] registers\[59\]\[37\]
+ _06301_ _06091_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__mux4_1
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18629_ registers\[12\]\[7\] registers\[13\]\[7\] registers\[14\]\[7\] registers\[15\]\[7\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__mux4_1
X_30907_ registers\[10\]\[17\] _12970_ _13933_ VGND VGND VPWR VPWR _13941_ sky130_fd_sc_hd__mux2_1
XFILLER_80_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34675_ clknet_leaf_408_CLK _02789_ VGND VGND VPWR VPWR registers\[26\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31887_ _14456_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21640_ registers\[16\]\[27\] registers\[17\]\[27\] registers\[18\]\[27\] registers\[19\]\[27\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__mux4_1
X_33626_ clknet_leaf_32_CLK _01740_ VGND VGND VPWR VPWR registers\[42\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_30838_ _13904_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33557_ clknet_leaf_125_CLK _01671_ VGND VGND VPWR VPWR registers\[43\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_21571_ _08075_ _08243_ _08244_ _08078_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__a22o_1
XFILLER_123_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30769_ _13868_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_11 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_22 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23310_ net48 VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__buf_4
X_20522_ registers\[56\]\[62\] registers\[57\]\[62\] registers\[58\]\[62\] registers\[59\]\[62\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__mux4_1
XANTENNA_33 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32508_ clknet_leaf_289_CLK _00622_ VGND VGND VPWR VPWR registers\[60\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_44 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ registers\[57\]\[14\] _10334_ _10326_ VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__mux2_1
X_33488_ clknet_leaf_129_CLK _01602_ VGND VGND VPWR VPWR registers\[44\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_55 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_66 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_77 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23241_ net25 VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__buf_4
X_35227_ clknet_leaf_6_CLK _03341_ VGND VGND VPWR VPWR registers\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_20453_ _07135_ _07142_ _07149_ _07156_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__or4_1
XANTENNA_88 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32439_ clknet_leaf_426_CLK _00553_ VGND VGND VPWR VPWR registers\[29\]\[41\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_99 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23172_ _09715_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
X_35158_ clknet_leaf_89_CLK _03272_ VGND VGND VPWR VPWR registers\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_20384_ _05060_ _07088_ _07089_ _05066_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__a22o_1
XFILLER_107_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34109_ clknet_leaf_276_CLK _02223_ VGND VGND VPWR VPWR registers\[35\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22123_ _08469_ _08779_ _08780_ _08472_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__a22o_1
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35089_ clknet_leaf_106_CLK _03203_ VGND VGND VPWR VPWR registers\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_27980_ _11740_ registers\[31\]\[5\] _12364_ VGND VGND VPWR VPWR _12370_ sky130_fd_sc_hd__mux2_1
Xoutput140 net140 VGND VGND VPWR VPWR D1[55] sky130_fd_sc_hd__buf_2
XTAP_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 net151 VGND VGND VPWR VPWR D1[7] sky130_fd_sc_hd__buf_2
XTAP_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput162 net162 VGND VGND VPWR VPWR D2[17] sky130_fd_sc_hd__buf_2
XFILLER_47_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 net173 VGND VGND VPWR VPWR D2[27] sky130_fd_sc_hd__buf_2
X_26931_ net29 VGND VGND VPWR VPWR _11803_ sky130_fd_sc_hd__clkbuf_4
X_22054_ registers\[52\]\[39\] registers\[53\]\[39\] registers\[54\]\[39\] registers\[55\]\[39\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__mux4_1
XTAP_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput184 net184 VGND VGND VPWR VPWR D2[37] sky130_fd_sc_hd__buf_2
XFILLER_216_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput195 net195 VGND VGND VPWR VPWR D2[47] sky130_fd_sc_hd__buf_2
XTAP_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ registers\[24\]\[9\] registers\[25\]\[9\] registers\[26\]\[9\] registers\[27\]\[9\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__mux4_1
XFILLER_247_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29650_ registers\[20\]\[62\] _13064_ _13210_ VGND VGND VPWR VPWR _13279_ sky130_fd_sc_hd__mux2_1
XFILLER_216_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26862_ _11756_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28601_ _12696_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25813_ _11197_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
X_26793_ registers\[40\]\[50\] _10409_ _11713_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__mux2_1
X_29581_ registers\[20\]\[29\] _12995_ _13233_ VGND VGND VPWR VPWR _13243_ sky130_fd_sc_hd__mux2_1
XFILLER_214_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25744_ _11161_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
X_28532_ _12660_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__clkbuf_1
X_22956_ _09566_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21907_ registers\[48\]\[35\] registers\[49\]\[35\] registers\[50\]\[35\] registers\[51\]\[35\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__mux4_1
X_28463_ _11818_ registers\[28\]\[42\] _12621_ VGND VGND VPWR VPWR _12624_ sky130_fd_sc_hd__mux2_1
X_25675_ registers\[48\]\[34\] _10376_ _11119_ VGND VGND VPWR VPWR _11124_ sky130_fd_sc_hd__mux2_1
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22887_ _09519_ registers\[62\]\[2\] _09515_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__mux2_1
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27414_ registers\[36\]\[58\] _10426_ _12062_ VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__mux2_1
X_24626_ _09556_ registers\[55\]\[20\] _10536_ VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__mux2_1
X_28394_ _12587_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__clkbuf_1
X_21838_ _08469_ _08502_ _08503_ _08472_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__a22o_1
XFILLER_197_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27345_ registers\[36\]\[25\] _10357_ _12029_ VGND VGND VPWR VPWR _12035_ sky130_fd_sc_hd__mux2_1
XFILLER_197_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24557_ _09626_ registers\[56\]\[53\] _10495_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__mux2_1
XFILLER_168_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21769_ registers\[36\]\[31\] registers\[37\]\[31\] registers\[38\]\[31\] registers\[39\]\[31\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__mux4_1
XFILLER_15_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23508_ _09912_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__clkbuf_1
X_27276_ _11998_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24488_ _09556_ registers\[56\]\[20\] _10462_ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__mux2_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29015_ registers\[24\]\[48\] _10405_ _12905_ VGND VGND VPWR VPWR _12914_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26227_ _10812_ registers\[44\]\[39\] _11405_ VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__mux2_1
X_23439_ _09876_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26158_ _10743_ registers\[44\]\[6\] _11372_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__mux2_1
XFILLER_164_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25109_ net32 VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__buf_2
XFILLER_180_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18980_ registers\[0\]\[17\] registers\[1\]\[17\] registers\[2\]\[17\] registers\[3\]\[17\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__mux4_1
X_26089_ _11342_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29917_ _13419_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__clkbuf_1
X_17931_ _14576_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__buf_6
XFILLER_124_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17862_ _14530_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__buf_4
X_29848_ _13383_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19601_ _06226_ _06327_ _06328_ _06231_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__a22o_1
X_16813_ registers\[32\]\[21\] registers\[33\]\[21\] registers\[34\]\[21\] registers\[35\]\[21\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15306_ sky130_fd_sc_hd__mux4_1
X_29779_ registers\[1\]\[59\] _13058_ _13337_ VGND VGND VPWR VPWR _13347_ sky130_fd_sc_hd__mux2_1
X_17793_ _04571_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31810_ _14415_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19532_ _06262_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__buf_2
XFILLER_235_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16744_ registers\[56\]\[19\] registers\[57\]\[19\] registers\[58\]\[19\] registers\[59\]\[19\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15239_ sky130_fd_sc_hd__mux4_1
X_32790_ clknet_leaf_65_CLK _00904_ VGND VGND VPWR VPWR registers\[55\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19463_ _06162_ _06171_ _06181_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__or4_1
X_31741_ _14379_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16675_ registers\[60\]\[17\] registers\[61\]\[17\] registers\[62\]\[17\] registers\[63\]\[17\]
+ _15070_ _14864_ VGND VGND VPWR VPWR _15172_ sky130_fd_sc_hd__mux4_1
XFILLER_235_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18414_ registers\[48\]\[1\] registers\[49\]\[1\] registers\[50\]\[1\] registers\[51\]\[1\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__mux4_1
XFILLER_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34460_ clknet_leaf_10_CLK _02574_ VGND VGND VPWR VPWR registers\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31672_ registers\[63\]\[60\] net57 _14276_ VGND VGND VPWR VPWR _14343_ sky130_fd_sc_hd__mux2_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ registers\[36\]\[29\] registers\[37\]\[29\] registers\[38\]\[29\] registers\[39\]\[29\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__mux4_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33411_ clknet_leaf_255_CLK _01525_ VGND VGND VPWR VPWR registers\[46\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_18345_ _05051_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__buf_8
X_30623_ registers\[12\]\[10\] _12955_ _13791_ VGND VGND VPWR VPWR _13792_ sky130_fd_sc_hd__mux2_1
X_34391_ clknet_leaf_98_CLK _02505_ VGND VGND VPWR VPWR registers\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36130_ clknet_leaf_46_CLK _04244_ VGND VGND VPWR VPWR registers\[49\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33342_ clknet_leaf_273_CLK _01456_ VGND VGND VPWR VPWR registers\[47\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18276_ _05038_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__buf_12
X_30554_ _13755_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput20 DW[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_4
X_17227_ registers\[28\]\[32\] registers\[29\]\[32\] registers\[30\]\[32\] registers\[31\]\[32\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15709_ sky130_fd_sc_hd__mux4_1
X_36061_ clknet_leaf_49_CLK _04175_ VGND VGND VPWR VPWR registers\[59\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33273_ clknet_leaf_337_CLK _01387_ VGND VGND VPWR VPWR registers\[48\]\[43\] sky130_fd_sc_hd__dfxtp_1
Xinput31 DW[37] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
XFILLER_239_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30485_ _09676_ registers\[13\]\[9\] _13709_ VGND VGND VPWR VPWR _13719_ sky130_fd_sc_hd__mux2_1
Xinput42 DW[47] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_6
X_35012_ clknet_leaf_202_CLK _03126_ VGND VGND VPWR VPWR registers\[21\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput53 DW[57] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_16
X_32224_ clknet_leaf_214_CLK _00338_ VGND VGND VPWR VPWR registers\[9\]\[55\] sky130_fd_sc_hd__dfxtp_1
Xinput64 DW[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_6
Xinput75 R2[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
XFILLER_200_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17158_ registers\[20\]\[30\] registers\[21\]\[30\] registers\[22\]\[30\] registers\[23\]\[30\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15642_ sky130_fd_sc_hd__mux4_1
Xinput86 RW[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16109_ _14573_ VGND VGND VPWR VPWR _14622_ sky130_fd_sc_hd__buf_4
XFILLER_157_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17089_ _14518_ VGND VGND VPWR VPWR _15574_ sky130_fd_sc_hd__buf_6
X_32155_ clknet_leaf_24_CLK _00269_ VGND VGND VPWR VPWR registers\[39\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31106_ _14045_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32086_ clknet_leaf_490_CLK _00062_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1044 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35914_ clknet_leaf_158_CLK _04028_ VGND VGND VPWR VPWR registers\[7\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_31037_ _14009_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35845_ clknet_leaf_220_CLK _03959_ VGND VGND VPWR VPWR registers\[8\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22810_ registers\[20\]\[61\] registers\[21\]\[61\] registers\[22\]\[61\] registers\[23\]\[61\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__mux4_1
X_35776_ clknet_leaf_242_CLK _03890_ VGND VGND VPWR VPWR registers\[0\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23790_ _10063_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
X_32988_ clknet_leaf_52_CLK _01102_ VGND VGND VPWR VPWR registers\[52\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22741_ _07276_ _09379_ _09380_ _07286_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__a22o_1
X_34727_ clknet_leaf_449_CLK _02841_ VGND VGND VPWR VPWR registers\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_213_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31939_ _14483_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25460_ _09651_ _09649_ _09650_ VGND VGND VPWR VPWR _11007_ sky130_fd_sc_hd__or3_1
X_22672_ registers\[56\]\[57\] registers\[57\]\[57\] registers\[58\]\[57\] registers\[59\]\[57\]
+ _09223_ _09013_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__mux4_1
X_34658_ clknet_leaf_474_CLK _02772_ VGND VGND VPWR VPWR registers\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24411_ registers\[57\]\[53\] _10416_ _10410_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__mux2_1
XFILLER_241_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33609_ clknet_leaf_245_CLK _01723_ VGND VGND VPWR VPWR registers\[43\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_21623_ _08126_ _08291_ _08294_ _08129_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25391_ _10971_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__clkbuf_1
X_34589_ clknet_leaf_7_CLK _02703_ VGND VGND VPWR VPWR registers\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27130_ _11837_ registers\[38\]\[51\] _11920_ VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__mux2_1
XFILLER_178_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24342_ net25 VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__buf_4
XFILLER_240_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21554_ registers\[48\]\[25\] registers\[49\]\[25\] registers\[50\]\[25\] registers\[51\]\[25\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__mux4_1
XFILLER_139_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20505_ _07203_ _07206_ _05133_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__o21ba_1
XFILLER_222_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27061_ _11885_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_1
X_24273_ net64 VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__buf_4
X_21485_ _08126_ _08159_ _08160_ _08129_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__a22o_1
XFILLER_222_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26012_ _11302_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
X_23224_ registers\[9\]\[26\] _09744_ _09735_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__mux2_1
X_20436_ registers\[52\]\[59\] registers\[53\]\[59\] registers\[54\]\[59\] registers\[55\]\[59\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__mux4_1
XFILLER_147_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23155_ _09651_ _09649_ _09650_ VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__or3b_1
XTAP_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20367_ _06912_ _07071_ _07072_ _06917_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__a22o_1
XFILLER_122_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22106_ _08761_ _08762_ _08763_ _08764_ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__a22o_1
XTAP_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23086_ _09653_ _09656_ VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__nor2_8
X_27963_ _12360_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1109 _14564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20298_ _06868_ _07005_ _07006_ _06871_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__a22o_1
XTAP_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29702_ registers\[1\]\[22\] _12981_ _13304_ VGND VGND VPWR VPWR _13307_ sky130_fd_sc_hd__mux2_1
XTAP_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26914_ _11791_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__clkbuf_1
X_22037_ _08423_ _08696_ _08697_ _08428_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__a22o_1
XFILLER_103_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27894_ _12324_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__clkbuf_1
XTAP_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29633_ _13270_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__clkbuf_1
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26845_ _11744_ registers\[3\]\[7\] _11730_ VGND VGND VPWR VPWR _11745_ sky130_fd_sc_hd__mux2_1
XTAP_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29564_ _13234_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23988_ _10168_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__clkbuf_1
X_26776_ registers\[40\]\[42\] _10393_ _11702_ VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__mux2_1
XFILLER_91_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28515_ _12651_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25727_ registers\[48\]\[59\] _10428_ _11141_ VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__mux2_1
X_22939_ _09554_ registers\[62\]\[19\] _09536_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__mux2_1
X_29495_ _09802_ registers\[21\]\[52\] _13195_ VGND VGND VPWR VPWR _13198_ sky130_fd_sc_hd__mux2_1
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16460_ registers\[32\]\[11\] registers\[33\]\[11\] registers\[34\]\[11\] registers\[35\]\[11\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _14963_ sky130_fd_sc_hd__mux4_1
X_28446_ _11801_ registers\[28\]\[34\] _12610_ VGND VGND VPWR VPWR _12615_ sky130_fd_sc_hd__mux2_1
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25658_ registers\[48\]\[26\] _10359_ _11108_ VGND VGND VPWR VPWR _11115_ sky130_fd_sc_hd__mux2_1
XFILLER_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16391_ registers\[56\]\[9\] registers\[57\]\[9\] registers\[58\]\[9\] registers\[59\]\[9\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _14896_ sky130_fd_sc_hd__mux4_1
X_24609_ _09540_ registers\[55\]\[12\] _10525_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__mux2_1
XFILLER_58_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28377_ _11732_ registers\[28\]\[1\] _12577_ VGND VGND VPWR VPWR _12579_ sky130_fd_sc_hd__mux2_1
X_25589_ registers\[4\]\[59\] _10428_ _11067_ VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__mux2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18130_ _04683_ _04896_ _04897_ _04686_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__a22o_1
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27328_ registers\[36\]\[17\] _10340_ _12018_ VGND VGND VPWR VPWR _12026_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18061_ _04637_ _04830_ _04831_ _04642_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__a22o_1
X_27259_ _11989_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17012_ _15295_ _15498_ _15499_ _15300_ VGND VGND VPWR VPWR _15500_ sky130_fd_sc_hd__a22o_1
XFILLER_176_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30270_ _13605_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_180_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_180_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18963_ registers\[40\]\[17\] registers\[41\]\[17\] registers\[42\]\[17\] registers\[43\]\[17\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__mux4_1
XFILLER_26_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1610 _15074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1621 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17914_ registers\[56\]\[52\] registers\[57\]\[52\] registers\[58\]\[52\] registers\[59\]\[52\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__mux4_1
XANTENNA_1632 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33960_ clknet_leaf_435_CLK _02074_ VGND VGND VPWR VPWR registers\[37\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1643 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18894_ registers\[32\]\[15\] registers\[33\]\[15\] registers\[34\]\[15\] registers\[35\]\[15\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__mux4_1
XTAP_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1654 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1665 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32911_ clknet_leaf_175_CLK _01025_ VGND VGND VPWR VPWR registers\[53\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1676 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17845_ registers\[8\]\[50\] registers\[9\]\[50\] registers\[10\]\[50\] registers\[11\]\[50\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__mux4_1
XFILLER_227_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1687 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33891_ clknet_leaf_47_CLK _02005_ VGND VGND VPWR VPWR registers\[38\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1698 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35630_ clknet_leaf_391_CLK _03744_ VGND VGND VPWR VPWR registers\[11\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_32842_ clknet_leaf_162_CLK _00956_ VGND VGND VPWR VPWR registers\[55\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_17776_ registers\[8\]\[48\] registers\[9\]\[48\] registers\[10\]\[48\] registers\[11\]\[48\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__mux4_1
XFILLER_94_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19515_ registers\[8\]\[32\] registers\[9\]\[32\] registers\[10\]\[32\] registers\[11\]\[32\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux4_1
X_35561_ clknet_leaf_398_CLK _03675_ VGND VGND VPWR VPWR registers\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_16727_ registers\[16\]\[18\] registers\[17\]\[18\] registers\[18\]\[18\] registers\[19\]\[18\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15223_ sky130_fd_sc_hd__mux4_1
XFILLER_35_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32773_ clknet_leaf_264_CLK _00887_ VGND VGND VPWR VPWR registers\[56\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_34512_ clknet_leaf_116_CLK _02626_ VGND VGND VPWR VPWR registers\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19446_ _06036_ _06177_ _06178_ _06039_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a22o_1
X_31724_ registers\[59\]\[20\] net13 _14370_ VGND VGND VPWR VPWR _14371_ sky130_fd_sc_hd__mux2_1
X_16658_ registers\[20\]\[16\] registers\[21\]\[16\] registers\[22\]\[16\] registers\[23\]\[16\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15156_ sky130_fd_sc_hd__mux4_1
X_35492_ clknet_leaf_467_CLK _03606_ VGND VGND VPWR VPWR registers\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34443_ clknet_leaf_150_CLK _02557_ VGND VGND VPWR VPWR registers\[30\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_31655_ _14334_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__clkbuf_1
X_19377_ _06036_ _06108_ _06111_ _06039_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__a22o_1
X_16589_ _14952_ _15087_ _15088_ _14957_ VGND VGND VPWR VPWR _15089_ sky130_fd_sc_hd__a22o_1
XFILLER_245_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30606_ registers\[12\]\[2\] _12939_ _13780_ VGND VGND VPWR VPWR _13783_ sky130_fd_sc_hd__mux2_1
XFILLER_176_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18328_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__buf_6
XFILLER_33_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34374_ clknet_leaf_213_CLK _02488_ VGND VGND VPWR VPWR registers\[31\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31586_ registers\[63\]\[19\] net11 _14288_ VGND VGND VPWR VPWR _14298_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_36__f_CLK clknet_5_18_0_CLK VGND VGND VPWR VPWR clknet_6_36__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_36113_ clknet_leaf_74_CLK _04227_ VGND VGND VPWR VPWR registers\[49\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33325_ clknet_leaf_344_CLK _01439_ VGND VGND VPWR VPWR registers\[47\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_18259_ registers\[8\]\[63\] registers\[9\]\[63\] registers\[10\]\[63\] registers\[11\]\[63\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux4_1
X_30537_ _13746_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36044_ clknet_leaf_167_CLK _04158_ VGND VGND VPWR VPWR registers\[63\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33256_ clknet_leaf_424_CLK _01370_ VGND VGND VPWR VPWR registers\[48\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_21270_ _07783_ _07948_ _07951_ _07786_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__a22o_1
X_30468_ _13710_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20221_ registers\[8\]\[52\] registers\[9\]\[52\] registers\[10\]\[52\] registers\[11\]\[52\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__mux4_1
X_32207_ clknet_leaf_353_CLK _00321_ VGND VGND VPWR VPWR registers\[9\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_171_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_171_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33187_ clknet_leaf_471_CLK _01301_ VGND VGND VPWR VPWR registers\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_30399_ _09758_ registers\[14\]\[32\] _13671_ VGND VGND VPWR VPWR _13674_ sky130_fd_sc_hd__mux2_1
XFILLER_172_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20152_ _06722_ _06863_ _06864_ _06725_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__a22o_1
XFILLER_172_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32138_ clknet_leaf_460_CLK _00056_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24960_ _10657_ VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__buf_4
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32069_ clknet_leaf_199_CLK _00247_ VGND VGND VPWR VPWR registers\[62\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_20083_ _06722_ _06794_ _06797_ _06725_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__a22o_1
XFILLER_135_1251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _10127_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24891_ _09550_ registers\[53\]\[17\] _10669_ VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__mux2_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23842_ _10091_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
X_26630_ _11627_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__clkbuf_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35828_ clknet_leaf_324_CLK _03942_ VGND VGND VPWR VPWR registers\[8\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_507 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26561_ _11591_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__clkbuf_1
X_35759_ clknet_leaf_378_CLK _03873_ VGND VGND VPWR VPWR registers\[0\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_23773_ _10054_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_518 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20985_ registers\[32\]\[9\] registers\[33\]\[9\] registers\[34\]\[9\] registers\[35\]\[9\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__mux4_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_529 _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28300_ registers\[2\]\[29\] _10365_ _12528_ VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__mux2_1
XFILLER_92_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22724_ _09364_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25512_ registers\[4\]\[22\] _10351_ _11034_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__mux2_1
X_29280_ _09687_ registers\[22\]\[14\] _13080_ VGND VGND VPWR VPWR _13085_ sky130_fd_sc_hd__mux2_1
X_26492_ _11554_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28231_ _12501_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__clkbuf_1
X_25443_ _10998_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22655_ _09294_ _09297_ _09102_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__o21ba_1
XFILLER_201_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21606_ _07377_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__buf_4
XFILLER_181_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28162_ _12465_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__clkbuf_1
X_25374_ _10962_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__clkbuf_1
X_22586_ _09226_ _09230_ _09091_ _09092_ VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__o211a_1
XFILLER_178_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27113_ _11820_ registers\[38\]\[43\] _11909_ VGND VGND VPWR VPWR _11913_ sky130_fd_sc_hd__mux2_1
X_24325_ _10358_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
X_28093_ _11853_ registers\[31\]\[59\] _12419_ VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__mux2_1
X_21537_ registers\[24\]\[24\] registers\[25\]\[24\] registers\[26\]\[24\] registers\[27\]\[24\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__mux4_1
XFILLER_154_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27044_ _11750_ registers\[38\]\[10\] _11876_ VGND VGND VPWR VPWR _11877_ sky130_fd_sc_hd__mux2_1
X_24256_ registers\[57\]\[3\] _10311_ _10305_ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__mux2_1
X_21468_ _08141_ _08144_ _08073_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__o21ba_1
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23207_ _09734_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
X_20419_ registers\[28\]\[58\] registers\[29\]\[58\] registers\[30\]\[58\] registers\[31\]\[58\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__mux4_1
XFILLER_134_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_162_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_162_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24187_ _10273_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21399_ _07382_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23138_ _09692_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
XTAP_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28995_ _12903_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__clkbuf_1
XTAP_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27946_ registers\[32\]\[53\] _10416_ _12348_ VGND VGND VPWR VPWR _12352_ sky130_fd_sc_hd__mux2_1
XTAP_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23069_ _09642_ registers\[62\]\[61\] _09514_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__mux2_1
XTAP_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27877_ registers\[32\]\[20\] _10346_ _12315_ VGND VGND VPWR VPWR _12316_ sky130_fd_sc_hd__mux2_1
XTAP_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29616_ _13261_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__clkbuf_1
X_17630_ registers\[60\]\[44\] registers\[61\]\[44\] registers\[62\]\[44\] registers\[63\]\[44\]
+ _04412_ _15893_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__mux4_1
X_26828_ _11733_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_1
XTAP_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17561_ registers\[56\]\[42\] registers\[57\]\[42\] registers\[58\]\[42\] registers\[59\]\[42\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__mux4_1
X_29547_ _13225_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26759_ registers\[40\]\[34\] _10376_ _11691_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19300_ registers\[12\]\[26\] registers\[13\]\[26\] registers\[14\]\[26\] registers\[15\]\[26\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__mux4_1
XFILLER_229_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16512_ registers\[12\]\[12\] registers\[13\]\[12\] registers\[14\]\[12\] registers\[15\]\[12\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _15014_ sky130_fd_sc_hd__mux4_1
XFILLER_232_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29478_ _09784_ registers\[21\]\[44\] _13184_ VGND VGND VPWR VPWR _13189_ sky130_fd_sc_hd__mux2_1
X_17492_ registers\[8\]\[40\] registers\[9\]\[40\] registers\[10\]\[40\] registers\[11\]\[40\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15966_ sky130_fd_sc_hd__mux4_1
XFILLER_225_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19231_ registers\[12\]\[24\] registers\[13\]\[24\] registers\[14\]\[24\] registers\[15\]\[24\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__mux4_1
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28429_ _11784_ registers\[28\]\[26\] _12599_ VGND VGND VPWR VPWR _12606_ sky130_fd_sc_hd__mux2_1
X_16443_ _14587_ VGND VGND VPWR VPWR _14947_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19162_ registers\[8\]\[22\] registers\[9\]\[22\] registers\[10\]\[22\] registers\[11\]\[22\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__mux4_1
X_31440_ _14221_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16374_ registers\[16\]\[8\] registers\[17\]\[8\] registers\[18\]\[8\] registers\[19\]\[8\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14880_ sky130_fd_sc_hd__mux4_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18113_ registers\[4\]\[58\] registers\[5\]\[58\] registers\[6\]\[58\] registers\[7\]\[58\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__mux4_1
XFILLER_129_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31371_ registers\[7\]\[45\] net40 _14179_ VGND VGND VPWR VPWR _14185_ sky130_fd_sc_hd__mux2_1
X_19093_ _05693_ _05834_ _05835_ _05696_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a22o_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33110_ clknet_leaf_68_CLK _01224_ VGND VGND VPWR VPWR registers\[50\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30322_ _13632_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__clkbuf_1
X_18044_ _04540_ _04813_ _04814_ _04546_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__a22o_1
XFILLER_173_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34090_ clknet_leaf_435_CLK _02204_ VGND VGND VPWR VPWR registers\[35\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33041_ clknet_leaf_74_CLK _01155_ VGND VGND VPWR VPWR registers\[51\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_153_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_153_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30253_ _13596_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30184_ registers\[16\]\[59\] _13058_ _13550_ VGND VGND VPWR VPWR _13560_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19995_ _05095_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__buf_4
XFILLER_141_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18946_ _05059_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__clkbuf_4
X_34992_ clknet_leaf_385_CLK _03106_ VGND VGND VPWR VPWR registers\[21\]\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1440 _05059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1451 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33943_ clknet_leaf_117_CLK _02057_ VGND VGND VPWR VPWR registers\[37\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1462 _05156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1473 _05328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18877_ _05345_ _05624_ _05625_ _05348_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a22o_1
XFILLER_239_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1484 _06807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1495 _07324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17828_ _04333_ _04603_ _04604_ _04338_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a22o_1
X_33874_ clknet_leaf_120_CLK _01988_ VGND VGND VPWR VPWR registers\[38\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35613_ clknet_leaf_486_CLK _03727_ VGND VGND VPWR VPWR registers\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32825_ clknet_leaf_287_CLK _00939_ VGND VGND VPWR VPWR registers\[55\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17759_ _04340_ _04536_ _04537_ _04343_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a22o_1
XFILLER_35_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35544_ clknet_leaf_475_CLK _03658_ VGND VGND VPWR VPWR registers\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_20770_ _07386_ _07465_ _07466_ _07396_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__a22o_1
X_32756_ clknet_leaf_350_CLK _00870_ VGND VGND VPWR VPWR registers\[56\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31707_ registers\[59\]\[12\] net4 _14359_ VGND VGND VPWR VPWR _14362_ sky130_fd_sc_hd__mux2_1
XFILLER_126_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19429_ _06155_ _06160_ _06161_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__o21ba_2
XFILLER_223_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35475_ clknet_leaf_77_CLK _03589_ VGND VGND VPWR VPWR registers\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32687_ clknet_leaf_367_CLK _00801_ VGND VGND VPWR VPWR registers\[57\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22440_ registers\[52\]\[50\] registers\[53\]\[50\] registers\[54\]\[50\] registers\[55\]\[50\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__mux4_1
X_34426_ clknet_leaf_184_CLK _02540_ VGND VGND VPWR VPWR registers\[30\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31638_ _14325_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22371_ registers\[60\]\[48\] registers\[61\]\[48\] registers\[62\]\[48\] registers\[63\]\[48\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__mux4_1
X_34357_ clknet_leaf_416_CLK _02471_ VGND VGND VPWR VPWR registers\[31\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31569_ _14289_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_392_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_392_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_191_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24110_ _10232_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__buf_4
X_33308_ clknet_leaf_29_CLK _01422_ VGND VGND VPWR VPWR registers\[47\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_21322_ _07363_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__buf_4
X_25090_ _10797_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34288_ clknet_leaf_348_CLK _02402_ VGND VGND VPWR VPWR registers\[32\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36027_ clknet_leaf_288_CLK _04141_ VGND VGND VPWR VPWR registers\[63\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_24041_ _10196_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_144_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_144_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33239_ clknet_leaf_69_CLK _01353_ VGND VGND VPWR VPWR registers\[48\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_21253_ _07377_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__buf_6
XFILLER_176_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20204_ registers\[40\]\[52\] registers\[41\]\[52\] registers\[42\]\[52\] registers\[43\]\[52\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux4_1
XFILLER_176_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21184_ registers\[24\]\[14\] registers\[25\]\[14\] registers\[26\]\[14\] registers\[27\]\[14\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__mux4_1
XFILLER_85_1267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27800_ registers\[33\]\[48\] _10405_ _12266_ VGND VGND VPWR VPWR _12275_ sky130_fd_sc_hd__mux2_1
X_20135_ _06841_ _06846_ _06847_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__o21ba_1
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28780_ _11728_ registers\[25\]\[0\] _12790_ VGND VGND VPWR VPWR _12791_ sky130_fd_sc_hd__mux2_1
X_25992_ _11291_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27731_ registers\[33\]\[15\] _10336_ _12233_ VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__mux2_1
X_20066_ registers\[48\]\[48\] registers\[49\]\[48\] registers\[50\]\[48\] registers\[51\]\[48\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux4_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24943_ _10704_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27662_ _12202_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__clkbuf_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24874_ _09533_ registers\[53\]\[9\] _10658_ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__mux2_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29401_ _13148_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__clkbuf_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26613_ _11618_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__clkbuf_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23825_ _10081_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_304 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27593_ _12166_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__clkbuf_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_337 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29332_ _09773_ registers\[22\]\[39\] _13102_ VGND VGND VPWR VPWR _13112_ sky130_fd_sc_hd__mux2_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26544_ _11581_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_348 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23756_ _10045_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_359 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20968_ _07361_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__buf_6
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22707_ _07385_ _09346_ _09347_ _07395_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__a22o_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29263_ _09670_ registers\[22\]\[6\] _13069_ VGND VGND VPWR VPWR _13076_ sky130_fd_sc_hd__mux2_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23687_ _10007_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26475_ _11545_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20899_ registers\[24\]\[6\] registers\[25\]\[6\] registers\[26\]\[6\] registers\[27\]\[6\]
+ _07524_ _07525_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__mux4_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28214_ _11839_ registers\[30\]\[52\] _12490_ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22638_ registers\[44\]\[56\] registers\[45\]\[56\] registers\[46\]\[56\] registers\[47\]\[56\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__mux4_1
X_25426_ _10989_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29194_ net41 VGND VGND VPWR VPWR _13031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25357_ _10953_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_1
X_28145_ _12456_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__clkbuf_1
X_22569_ _09191_ _09198_ _09207_ _09214_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_383_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_383_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16090_ _14603_ VGND VGND VPWR VPWR _14604_ sky130_fd_sc_hd__buf_4
X_24308_ _10304_ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__buf_4
X_28076_ _12420_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25288_ _10916_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27027_ _11734_ registers\[38\]\[2\] _11865_ VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__mux2_1
X_24239_ _10300_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_135_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_135_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18800_ _05547_ _05548_ _05549_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__a22o_1
XFILLER_123_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19780_ _06233_ _06501_ _06502_ _06236_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__a22o_1
XFILLER_231_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28978_ registers\[24\]\[30\] _10367_ _12894_ VGND VGND VPWR VPWR _12895_ sky130_fd_sc_hd__mux2_1
X_16992_ _15206_ _15476_ _15479_ _15210_ VGND VGND VPWR VPWR _15480_ sky130_fd_sc_hd__a22o_1
XFILLER_235_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18731_ _05104_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__buf_4
XTAP_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27929_ registers\[32\]\[45\] _10399_ _12337_ VGND VGND VPWR VPWR _12343_ sky130_fd_sc_hd__mux2_1
XTAP_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _05412_ _05414_ _05415_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__a22o_1
XFILLER_7_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30940_ _13958_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_237_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17613_ registers\[20\]\[43\] registers\[21\]\[43\] registers\[22\]\[43\] registers\[23\]\[43\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__mux4_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30871_ _13921_ VGND VGND VPWR VPWR _13922_ sky130_fd_sc_hd__buf_4
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18593_ _05059_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__buf_4
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32610_ clknet_leaf_45_CLK _00724_ VGND VGND VPWR VPWR registers\[58\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_17544_ _04294_ _04328_ _04329_ _04299_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a22o_1
XFILLER_45_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33590_ clknet_leaf_341_CLK _01704_ VGND VGND VPWR VPWR registers\[43\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_860 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_871 _09509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32541_ clknet_leaf_473_CLK _00655_ VGND VGND VPWR VPWR registers\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_882 _09554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17475_ _15677_ _15947_ _15948_ _15682_ VGND VGND VPWR VPWR _15949_ sky130_fd_sc_hd__a22o_1
XANTENNA_893 _09648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19214_ _05883_ _05951_ _05952_ _05888_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__a22o_1
X_35260_ clknet_leaf_190_CLK _03374_ VGND VGND VPWR VPWR registers\[17\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16426_ _14855_ _14928_ _14929_ _14861_ VGND VGND VPWR VPWR _14930_ sky130_fd_sc_hd__a22o_1
XFILLER_73_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32472_ clknet_leaf_54_CLK _00586_ VGND VGND VPWR VPWR registers\[60\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34211_ clknet_leaf_56_CLK _02325_ VGND VGND VPWR VPWR registers\[33\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31423_ _14212_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__clkbuf_1
X_19145_ registers\[40\]\[22\] registers\[41\]\[22\] registers\[42\]\[22\] registers\[43\]\[22\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__mux4_1
X_16357_ _14539_ VGND VGND VPWR VPWR _14863_ sky130_fd_sc_hd__clkbuf_4
X_35191_ clknet_leaf_310_CLK _03305_ VGND VGND VPWR VPWR registers\[18\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_374_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_374_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34142_ clknet_leaf_22_CLK _02256_ VGND VGND VPWR VPWR registers\[34\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31354_ registers\[7\]\[37\] net31 _14168_ VGND VGND VPWR VPWR _14176_ sky130_fd_sc_hd__mux2_1
X_19076_ _05812_ _05817_ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__o21ba_1
X_16288_ _14490_ VGND VGND VPWR VPWR _14796_ sky130_fd_sc_hd__buf_4
XFILLER_201_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_5_31_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_31_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_161_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18027_ registers\[16\]\[55\] registers\[17\]\[55\] registers\[18\]\[55\] registers\[19\]\[55\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux4_1
X_30305_ registers\[15\]\[52\] _13044_ _13621_ VGND VGND VPWR VPWR _13624_ sky130_fd_sc_hd__mux2_1
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_126_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_161_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34073_ clknet_leaf_91_CLK _02187_ VGND VGND VPWR VPWR registers\[35\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_31285_ registers\[7\]\[4\] net45 _14135_ VGND VGND VPWR VPWR _14140_ sky130_fd_sc_hd__mux2_1
X_33024_ clknet_leaf_267_CLK _01138_ VGND VGND VPWR VPWR registers\[52\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30236_ _13587_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30167_ _13551_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__clkbuf_1
X_19978_ registers\[28\]\[45\] registers\[29\]\[45\] registers\[30\]\[45\] registers\[31\]\[45\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__mux4_1
XFILLER_228_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ registers\[36\]\[16\] registers\[37\]\[16\] registers\[38\]\[16\] registers\[39\]\[16\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__mux4_1
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34975_ clknet_leaf_490_CLK _03089_ VGND VGND VPWR VPWR registers\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_30098_ registers\[16\]\[18\] _12972_ _13506_ VGND VGND VPWR VPWR _13515_ sky130_fd_sc_hd__mux2_1
XANTENNA_1270 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1281 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1292 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21940_ _08326_ _08601_ _08602_ _08332_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__a22o_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33926_ clknet_leaf_246_CLK _02040_ VGND VGND VPWR VPWR registers\[38\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33857_ clknet_leaf_240_CLK _01971_ VGND VGND VPWR VPWR registers\[3\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21871_ _08532_ _08535_ _08397_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__o21ba_1
XFILLER_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23610_ _09967_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
X_20822_ registers\[8\]\[4\] registers\[9\]\[4\] registers\[10\]\[4\] registers\[11\]\[4\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__mux4_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32808_ clknet_leaf_423_CLK _00922_ VGND VGND VPWR VPWR registers\[55\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24590_ _09521_ registers\[55\]\[3\] _10514_ VGND VGND VPWR VPWR _10518_ sky130_fd_sc_hd__mux2_1
X_33788_ clknet_leaf_277_CLK _01902_ VGND VGND VPWR VPWR registers\[40\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23541_ _09628_ registers\[19\]\[54\] _09925_ VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__mux2_1
X_35527_ clknet_leaf_214_CLK _03641_ VGND VGND VPWR VPWR registers\[13\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_20753_ registers\[52\]\[2\] registers\[53\]\[2\] registers\[54\]\[2\] registers\[55\]\[2\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__mux4_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32739_ clknet_leaf_443_CLK _00853_ VGND VGND VPWR VPWR registers\[56\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26260_ _11432_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35458_ clknet_leaf_239_CLK _03572_ VGND VGND VPWR VPWR registers\[14\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23472_ _09559_ registers\[19\]\[21\] _09892_ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__mux2_1
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20684_ _07382_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_206_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25211_ _10864_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__buf_4
X_22423_ _09069_ _09072_ _08773_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__o21ba_1
X_34409_ clknet_leaf_404_CLK _02523_ VGND VGND VPWR VPWR registers\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26191_ _11396_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
X_35389_ clknet_leaf_298_CLK _03503_ VGND VGND VPWR VPWR registers\[15\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_365_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_365_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25142_ _10832_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__clkbuf_1
X_22354_ registers\[40\]\[48\] registers\[41\]\[48\] registers\[42\]\[48\] registers\[43\]\[48\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__mux4_1
XFILLER_104_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21305_ _07278_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_117_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_117_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_29950_ _13437_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__clkbuf_1
X_25073_ _10785_ registers\[52\]\[26\] _10773_ VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__mux2_1
XFILLER_219_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22285_ registers\[32\]\[46\] registers\[33\]\[46\] registers\[34\]\[46\] registers\[35\]\[46\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__mux4_1
XFILLER_3_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28901_ _11851_ registers\[25\]\[58\] _12845_ VGND VGND VPWR VPWR _12854_ sky130_fd_sc_hd__mux2_1
X_24024_ _10187_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21236_ _07331_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__buf_4
XFILLER_172_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29881_ registers\[18\]\[43\] _13025_ _13397_ VGND VGND VPWR VPWR _13401_ sky130_fd_sc_hd__mux2_1
XFILLER_236_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28832_ _11782_ registers\[25\]\[25\] _12812_ VGND VGND VPWR VPWR _12818_ sky130_fd_sc_hd__mux2_1
X_21167_ registers\[56\]\[14\] registers\[57\]\[14\] registers\[58\]\[14\] registers\[59\]\[14\]
+ _07851_ _07641_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20118_ registers\[16\]\[49\] registers\[17\]\[49\] registers\[18\]\[49\] registers\[19\]\[49\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__mux4_1
XFILLER_63_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28763_ _12781_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__clkbuf_1
X_25975_ _11282_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21098_ registers\[36\]\[12\] registers\[37\]\[12\] registers\[38\]\[12\] registers\[39\]\[12\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__mux4_1
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27714_ registers\[33\]\[7\] _10319_ _12222_ VGND VGND VPWR VPWR _12230_ sky130_fd_sc_hd__mux2_1
X_20049_ registers\[20\]\[47\] registers\[21\]\[47\] registers\[22\]\[47\] registers\[23\]\[47\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__mux4_1
X_24926_ _10695_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28694_ _12745_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27645_ _12193_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24857_ _10659_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_112 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_123 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_861 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23808_ _09619_ registers\[29\]\[50\] _10072_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__mux2_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27576_ _12157_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__clkbuf_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24788_ _09582_ registers\[54\]\[32\] _10620_ VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__mux2_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_156 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_167 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29315_ _13103_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__clkbuf_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26527_ _10842_ registers\[42\]\[53\] _11569_ VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__mux2_1
XANTENNA_178 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23739_ _10036_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_189 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29246_ net60 VGND VGND VPWR VPWR _13066_ sky130_fd_sc_hd__buf_2
XFILLER_186_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17260_ registers\[20\]\[33\] registers\[21\]\[33\] registers\[22\]\[33\] registers\[23\]\[33\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15741_ sky130_fd_sc_hd__mux4_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26458_ _10772_ registers\[42\]\[20\] _11536_ VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__mux2_1
XFILLER_109_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16211_ _14655_ _14719_ _14720_ _14658_ VGND VGND VPWR VPWR _14721_ sky130_fd_sc_hd__a22o_1
XFILLER_201_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25409_ _10980_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__clkbuf_1
X_29177_ registers\[23\]\[40\] _13018_ _13019_ VGND VGND VPWR VPWR _13020_ sky130_fd_sc_hd__mux2_1
X_17191_ _15638_ _15672_ _15673_ _15643_ VGND VGND VPWR VPWR _15674_ sky130_fd_sc_hd__a22o_1
XFILLER_35_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_356_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_356_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_224_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26389_ _11500_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16142_ _14648_ _14651_ _14652_ _14653_ VGND VGND VPWR VPWR _14654_ sky130_fd_sc_hd__a22o_1
X_28128_ _11753_ registers\[30\]\[11\] _12446_ VGND VGND VPWR VPWR _12448_ sky130_fd_sc_hd__mux2_1
XFILLER_143_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_108_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16073_ _14489_ VGND VGND VPWR VPWR _14587_ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28059_ _12411_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19901_ registers\[0\]\[43\] registers\[1\]\[43\] registers\[2\]\[43\] registers\[3\]\[43\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__mux4_1
X_31070_ registers\[0\]\[30\] _12997_ _14026_ VGND VGND VPWR VPWR _14027_ sky130_fd_sc_hd__mux2_1
XFILLER_170_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30021_ _13474_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19832_ registers\[8\]\[41\] registers\[9\]\[41\] registers\[10\]\[41\] registers\[11\]\[41\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__mux4_1
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19763_ _06483_ _06486_ _06180_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__o21ba_1
X_16975_ _15460_ _15463_ _15302_ VGND VGND VPWR VPWR _15464_ sky130_fd_sc_hd__o21ba_1
X_18714_ registers\[40\]\[10\] registers\[41\]\[10\] registers\[42\]\[10\] registers\[43\]\[10\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__mux4_1
X_34760_ clknet_leaf_218_CLK _02874_ VGND VGND VPWR VPWR registers\[25\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31972_ clknet_leaf_5_CLK _00142_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_1
X_19694_ _06182_ _06418_ _06419_ _06185_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__a22o_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 DW[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_8
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33711_ clknet_leaf_360_CLK _01825_ VGND VGND VPWR VPWR registers\[41\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_18645_ registers\[44\]\[8\] registers\[45\]\[8\] registers\[46\]\[8\] registers\[47\]\[8\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__mux4_1
XFILLER_225_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30923_ _13949_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__clkbuf_1
X_34691_ clknet_leaf_223_CLK _02805_ VGND VGND VPWR VPWR registers\[26\]\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33642_ clknet_leaf_428_CLK _01756_ VGND VGND VPWR VPWR registers\[42\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_30854_ _09810_ registers\[11\]\[56\] _13906_ VGND VGND VPWR VPWR _13913_ sky130_fd_sc_hd__mux2_1
X_18576_ registers\[36\]\[6\] registers\[37\]\[6\] registers\[38\]\[6\] registers\[39\]\[6\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__mux4_1
XFILLER_36_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ _15884_ _04311_ _04312_ _15890_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__a22o_1
XFILLER_221_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33573_ clknet_leaf_57_CLK _01687_ VGND VGND VPWR VPWR registers\[43\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30785_ _09730_ registers\[11\]\[23\] _13873_ VGND VGND VPWR VPWR _13877_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_690 _06643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35312_ clknet_leaf_393_CLK _03426_ VGND VGND VPWR VPWR registers\[16\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32524_ clknet_leaf_167_CLK _00638_ VGND VGND VPWR VPWR registers\[60\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17458_ registers\[0\]\[39\] registers\[1\]\[39\] registers\[2\]\[39\] registers\[3\]\[39\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15933_ sky130_fd_sc_hd__mux4_1
XFILLER_178_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16409_ registers\[20\]\[9\] registers\[21\]\[9\] registers\[22\]\[9\] registers\[23\]\[9\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14914_ sky130_fd_sc_hd__mux4_1
X_35243_ clknet_leaf_408_CLK _03357_ VGND VGND VPWR VPWR registers\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_32455_ clknet_leaf_206_CLK _00569_ VGND VGND VPWR VPWR registers\[29\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_347_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_347_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17389_ registers\[4\]\[37\] registers\[5\]\[37\] registers\[6\]\[37\] registers\[7\]\[37\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15866_ sky130_fd_sc_hd__mux4_1
X_31406_ registers\[7\]\[62\] net59 _14134_ VGND VGND VPWR VPWR _14203_ sky130_fd_sc_hd__mux2_1
X_19128_ _05688_ _05868_ _05869_ _05691_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__a22o_1
XFILLER_192_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35174_ clknet_leaf_449_CLK _03288_ VGND VGND VPWR VPWR registers\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32386_ clknet_leaf_264_CLK _00500_ VGND VGND VPWR VPWR registers\[61\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34125_ clknet_leaf_170_CLK _02239_ VGND VGND VPWR VPWR registers\[35\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_31337_ registers\[7\]\[29\] net22 _14157_ VGND VGND VPWR VPWR _14167_ sky130_fd_sc_hd__mux2_1
X_19059_ registers\[16\]\[19\] registers\[17\]\[19\] registers\[18\]\[19\] registers\[19\]\[19\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__mux4_1
X_34056_ clknet_leaf_237_CLK _02170_ VGND VGND VPWR VPWR registers\[36\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_22070_ _08726_ _08729_ _08430_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__o21ba_1
X_31268_ _14130_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21021_ _07440_ _07708_ _07709_ _07443_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__a22o_1
X_33007_ clknet_leaf_368_CLK _01121_ VGND VGND VPWR VPWR registers\[52\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_30219_ registers\[15\]\[11\] _12958_ _13577_ VGND VGND VPWR VPWR _13579_ sky130_fd_sc_hd__mux2_1
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31199_ _14094_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25760_ _11169_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
X_22972_ net24 VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__clkbuf_4
X_34958_ clknet_leaf_115_CLK _03072_ VGND VGND VPWR VPWR registers\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24711_ _09642_ registers\[55\]\[61\] _10513_ VGND VGND VPWR VPWR _10581_ sky130_fd_sc_hd__mux2_1
XFILLER_56_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21923_ registers\[16\]\[35\] registers\[17\]\[35\] registers\[18\]\[35\] registers\[19\]\[35\]
+ _08279_ _08280_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__mux4_1
X_33909_ clknet_leaf_343_CLK _02023_ VGND VGND VPWR VPWR registers\[38\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25691_ _11132_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34889_ clknet_leaf_212_CLK _03003_ VGND VGND VPWR VPWR registers\[23\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_27430_ _11732_ registers\[35\]\[1\] _12078_ VGND VGND VPWR VPWR _12080_ sky130_fd_sc_hd__mux2_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _08272_ _08518_ _08519_ _08275_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__a22o_1
XFILLER_58_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24642_ _09573_ registers\[55\]\[28\] _10536_ VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__mux2_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20805_ _07500_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_2
XFILLER_169_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27361_ _12043_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__clkbuf_1
X_24573_ _09642_ registers\[56\]\[61\] _10439_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__mux2_1
XFILLER_24_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21785_ _08449_ _08452_ _08416_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__o21ba_1
XFILLER_230_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29100_ _12967_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__clkbuf_1
X_26312_ _10762_ registers\[43\]\[15\] _11454_ VGND VGND VPWR VPWR _11460_ sky130_fd_sc_hd__mux2_1
X_20736_ _07275_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__buf_4
XFILLER_195_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23524_ _09611_ registers\[19\]\[46\] _09914_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__mux2_1
X_27292_ _12006_ VGND VGND VPWR VPWR _12007_ sky130_fd_sc_hd__buf_4
XFILLER_93_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29031_ _12922_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26243_ _11423_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_1
X_23455_ _09542_ registers\[19\]\[13\] _09881_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__mux2_1
X_20667_ _07300_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_338_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_338_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22406_ registers\[60\]\[49\] registers\[61\]\[49\] registers\[62\]\[49\] registers\[63\]\[49\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__mux4_1
XFILLER_17_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23386_ registers\[39\]\[46\] _09788_ _09840_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__mux2_1
X_26174_ _11387_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20598_ _07287_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__buf_4
XFILLER_221_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22337_ _08985_ _08988_ _08748_ _08749_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__o211a_1
X_25125_ net38 VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__buf_2
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29933_ _13428_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__clkbuf_1
X_25056_ _10774_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
X_22268_ registers\[8\]\[45\] registers\[9\]\[45\] registers\[10\]\[45\] registers\[11\]\[45\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__mux4_1
XFILLER_65_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24007_ _10178_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
X_21219_ registers\[28\]\[15\] registers\[29\]\[15\] registers\[30\]\[15\] registers\[31\]\[15\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__mux4_1
X_29864_ registers\[18\]\[35\] _13008_ _13386_ VGND VGND VPWR VPWR _13392_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22199_ _08851_ _08854_ _08748_ _08749_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__o211a_1
XFILLER_239_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28815_ _11765_ registers\[25\]\[17\] _12801_ VGND VGND VPWR VPWR _12809_ sky130_fd_sc_hd__mux2_1
X_29795_ registers\[18\]\[2\] _12939_ _13353_ VGND VGND VPWR VPWR _13356_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28746_ _12772_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__clkbuf_1
X_16760_ _14947_ _15253_ _15254_ _14950_ VGND VGND VPWR VPWR _15255_ sky130_fd_sc_hd__a22o_1
XFILLER_59_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25958_ _11273_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
X_24909_ _10686_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
X_16691_ _14952_ _15186_ _15187_ _14957_ VGND VGND VPWR VPWR _15188_ sky130_fd_sc_hd__a22o_1
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28677_ _12736_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__clkbuf_1
X_25889_ _11237_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18430_ registers\[28\]\[1\] registers\[29\]\[1\] registers\[30\]\[1\] registers\[31\]\[1\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__mux4_1
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27628_ registers\[34\]\[30\] _10367_ _12184_ VGND VGND VPWR VPWR _12185_ sky130_fd_sc_hd__mux2_1
XFILLER_234_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ registers\[12\]\[0\] registers\[13\]\[0\] registers\[14\]\[0\] registers\[15\]\[0\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__mux4_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27559_ _11861_ registers\[35\]\[63\] _12077_ VGND VGND VPWR VPWR _12147_ sky130_fd_sc_hd__mux2_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _15787_ _15790_ _15620_ _15621_ VGND VGND VPWR VPWR _15791_ sky130_fd_sc_hd__o211a_1
XFILLER_30_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18292_ registers\[32\]\[0\] registers\[33\]\[0\] registers\[34\]\[0\] registers\[35\]\[0\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__mux4_1
XFILLER_226_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30570_ _13763_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__clkbuf_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29229_ registers\[23\]\[57\] _13054_ _13040_ VGND VGND VPWR VPWR _13055_ sky130_fd_sc_hd__mux2_1
X_17243_ registers\[60\]\[33\] registers\[61\]\[33\] registers\[62\]\[33\] registers\[63\]\[33\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15724_ sky130_fd_sc_hd__mux4_1
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_329_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_329_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32240_ clknet_leaf_365_CLK _00354_ VGND VGND VPWR VPWR registers\[39\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_17174_ _15541_ _15655_ _15656_ _15547_ VGND VGND VPWR VPWR _15657_ sky130_fd_sc_hd__a22o_1
XFILLER_31_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16125_ _14570_ _14636_ _14637_ _14582_ VGND VGND VPWR VPWR _14638_ sky130_fd_sc_hd__a22o_1
XFILLER_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32171_ clknet_leaf_440_CLK _00285_ VGND VGND VPWR VPWR registers\[39\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31122_ registers\[0\]\[55\] _13050_ _14048_ VGND VGND VPWR VPWR _14054_ sky130_fd_sc_hd__mux2_1
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16056_ _14510_ VGND VGND VPWR VPWR _14570_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31053_ registers\[0\]\[22\] _12981_ _14015_ VGND VGND VPWR VPWR _14018_ sky130_fd_sc_hd__mux2_1
X_35930_ clknet_leaf_476_CLK _04044_ VGND VGND VPWR VPWR registers\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30004_ _13465_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__clkbuf_1
X_19815_ _06529_ _06536_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__o21ba_1
X_35861_ clknet_leaf_78_CLK _03975_ VGND VGND VPWR VPWR registers\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34812_ clknet_leaf_306_CLK _02926_ VGND VGND VPWR VPWR registers\[24\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_16958_ _15206_ _15445_ _15446_ _15210_ VGND VGND VPWR VPWR _15447_ sky130_fd_sc_hd__a22o_1
X_19746_ registers\[44\]\[39\] registers\[45\]\[39\] registers\[46\]\[39\] registers\[47\]\[39\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__mux4_1
XFILLER_244_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35792_ clknet_leaf_136_CLK _03906_ VGND VGND VPWR VPWR registers\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31955_ clknet_leaf_0_CLK _00183_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
X_19677_ _06397_ _06402_ _06161_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21ba_1
X_34743_ clknet_leaf_426_CLK _02857_ VGND VGND VPWR VPWR registers\[25\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16889_ _15198_ _15378_ _15379_ _15204_ VGND VGND VPWR VPWR _15380_ sky130_fd_sc_hd__a22o_1
XFILLER_77_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18628_ _05345_ _05382_ _05383_ _05348_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__a22o_1
X_30906_ _13940_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__clkbuf_1
X_34674_ clknet_leaf_412_CLK _02788_ VGND VGND VPWR VPWR registers\[26\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31886_ _09760_ registers\[49\]\[33\] _14452_ VGND VGND VPWR VPWR _14456_ sky130_fd_sc_hd__mux2_1
XFILLER_212_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33625_ clknet_leaf_90_CLK _01739_ VGND VGND VPWR VPWR registers\[42\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_30837_ _09793_ registers\[11\]\[48\] _13895_ VGND VGND VPWR VPWR _13904_ sky130_fd_sc_hd__mux2_1
X_18559_ registers\[12\]\[5\] registers\[13\]\[5\] registers\[14\]\[5\] registers\[15\]\[5\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__mux4_1
XFILLER_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33556_ clknet_leaf_119_CLK _01670_ VGND VGND VPWR VPWR registers\[43\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_21570_ registers\[16\]\[25\] registers\[17\]\[25\] registers\[18\]\[25\] registers\[19\]\[25\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__mux4_1
X_30768_ _09689_ registers\[11\]\[15\] _13862_ VGND VGND VPWR VPWR _13868_ sky130_fd_sc_hd__mux2_1
XFILLER_33_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20521_ _07218_ _07221_ _05073_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__o21ba_1
X_32507_ clknet_leaf_288_CLK _00621_ VGND VGND VPWR VPWR registers\[60\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_23 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33487_ clknet_leaf_130_CLK _01601_ VGND VGND VPWR VPWR registers\[44\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30699_ _13831_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_45 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_56 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23240_ _09755_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
X_20452_ _07152_ _07155_ _06880_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__o21ba_1
XFILLER_119_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_78 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35226_ clknet_leaf_7_CLK _03340_ VGND VGND VPWR VPWR registers\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_32438_ clknet_leaf_419_CLK _00552_ VGND VGND VPWR VPWR registers\[29\]\[40\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_89 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23171_ registers\[9\]\[5\] _09668_ _09709_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__mux2_1
X_35157_ clknet_leaf_91_CLK _03271_ VGND VGND VPWR VPWR registers\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20383_ registers\[4\]\[57\] registers\[5\]\[57\] registers\[6\]\[57\] registers\[7\]\[57\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux4_1
X_32369_ clknet_leaf_371_CLK _00483_ VGND VGND VPWR VPWR registers\[61\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34108_ clknet_leaf_276_CLK _02222_ VGND VGND VPWR VPWR registers\[35\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_22122_ registers\[36\]\[41\] registers\[37\]\[41\] registers\[38\]\[41\] registers\[39\]\[41\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__mux4_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35088_ clknet_leaf_135_CLK _03202_ VGND VGND VPWR VPWR registers\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput130 net130 VGND VGND VPWR VPWR D1[46] sky130_fd_sc_hd__buf_2
XFILLER_115_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput141 net141 VGND VGND VPWR VPWR D1[56] sky130_fd_sc_hd__buf_2
XTAP_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput152 net152 VGND VGND VPWR VPWR D1[8] sky130_fd_sc_hd__buf_2
XTAP_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput163 net163 VGND VGND VPWR VPWR D2[18] sky130_fd_sc_hd__buf_2
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26930_ _11802_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_1
X_22053_ registers\[60\]\[39\] registers\[61\]\[39\] registers\[62\]\[39\] registers\[63\]\[39\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__mux4_1
X_34039_ clknet_leaf_340_CLK _02153_ VGND VGND VPWR VPWR registers\[36\]\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput174 net174 VGND VGND VPWR VPWR D2[28] sky130_fd_sc_hd__buf_2
XFILLER_115_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput185 net185 VGND VGND VPWR VPWR D2[38] sky130_fd_sc_hd__buf_2
Xoutput196 net196 VGND VGND VPWR VPWR D2[48] sky130_fd_sc_hd__buf_2
X_21004_ _07690_ _07693_ _07370_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__o21ba_1
XFILLER_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26861_ _11755_ registers\[3\]\[12\] _11751_ VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__mux2_1
XTAP_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28600_ _11820_ registers\[27\]\[43\] _12692_ VGND VGND VPWR VPWR _12696_ sky130_fd_sc_hd__mux2_1
XFILLER_60_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25812_ _10802_ registers\[47\]\[34\] _11192_ VGND VGND VPWR VPWR _11197_ sky130_fd_sc_hd__mux2_1
X_29580_ _13242_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__clkbuf_1
X_26792_ _11657_ VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__buf_4
XFILLER_112_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28531_ _11750_ registers\[27\]\[10\] _12659_ VGND VGND VPWR VPWR _12660_ sky130_fd_sc_hd__mux2_1
X_25743_ _10733_ registers\[47\]\[1\] _11159_ VGND VGND VPWR VPWR _11161_ sky130_fd_sc_hd__mux2_1
XFILLER_228_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22955_ _09565_ registers\[62\]\[24\] _09557_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__mux2_1
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21906_ registers\[56\]\[35\] registers\[57\]\[35\] registers\[58\]\[35\] registers\[59\]\[35\]
+ _08537_ _08327_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__mux4_1
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28462_ _12623_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25674_ _11123_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
X_22886_ net23 VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_216_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27413_ _12070_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24625_ _10513_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__buf_4
XFILLER_231_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28393_ _11748_ registers\[28\]\[9\] _12577_ VGND VGND VPWR VPWR _12587_ sky130_fd_sc_hd__mux2_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21837_ registers\[36\]\[33\] registers\[37\]\[33\] registers\[38\]\[33\] registers\[39\]\[33\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__mux4_1
XFILLER_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27344_ _12034_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__clkbuf_1
X_24556_ _10498_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21768_ registers\[44\]\[31\] registers\[45\]\[31\] registers\[46\]\[31\] registers\[47\]\[31\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__mux4_2
XFILLER_196_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20719_ _07413_ _07416_ _07339_ _07341_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__o211a_1
XFILLER_19_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23507_ _09594_ registers\[19\]\[38\] _09903_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27275_ _11847_ registers\[37\]\[56\] _11991_ VGND VGND VPWR VPWR _11998_ sky130_fd_sc_hd__mux2_1
XFILLER_200_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21699_ _08326_ _08367_ _08368_ _08332_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__a22o_1
X_24487_ _10439_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__buf_4
XFILLER_196_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29014_ _12913_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26226_ _11414_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
X_23438_ _09525_ registers\[19\]\[5\] _09870_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__mux2_1
XFILLER_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26157_ _11378_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
X_23369_ registers\[39\]\[38\] _09771_ _09829_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__mux2_1
XFILLER_152_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25108_ _10809_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26088_ _10808_ registers\[45\]\[37\] _11334_ VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__mux2_1
XFILLER_180_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17930_ _04632_ _04703_ _04704_ _04635_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a22o_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29916_ registers\[18\]\[60\] _13060_ _13352_ VGND VGND VPWR VPWR _13419_ sky130_fd_sc_hd__mux2_1
X_25039_ _10762_ registers\[52\]\[15\] _10752_ VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__mux2_1
XFILLER_117_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17861_ registers\[28\]\[50\] registers\[29\]\[50\] registers\[30\]\[50\] registers\[31\]\[50\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__mux4_1
XFILLER_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29847_ registers\[18\]\[27\] _12991_ _13375_ VGND VGND VPWR VPWR _13383_ sky130_fd_sc_hd__mux2_1
XFILLER_65_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19600_ registers\[32\]\[35\] registers\[33\]\[35\] registers\[34\]\[35\] registers\[35\]\[35\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__mux4_1
XFILLER_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16812_ registers\[40\]\[21\] registers\[41\]\[21\] registers\[42\]\[21\] registers\[43\]\[21\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15305_ sky130_fd_sc_hd__mux4_1
XFILLER_238_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29778_ _13346_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__clkbuf_1
X_17792_ _04539_ _04554_ _04563_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or4_2
XFILLER_226_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19531_ _06238_ _06245_ _06252_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__or4_1
X_28729_ _11813_ registers\[26\]\[40\] _12763_ VGND VGND VPWR VPWR _12764_ sky130_fd_sc_hd__mux2_1
X_16743_ _15234_ _15237_ _14926_ VGND VGND VPWR VPWR _15238_ sky130_fd_sc_hd__o21ba_1
XFILLER_98_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19462_ _06186_ _06193_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__o21ba_1
X_31740_ registers\[59\]\[28\] net21 _14370_ VGND VGND VPWR VPWR _14379_ sky130_fd_sc_hd__mux2_1
XFILLER_228_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16674_ _14855_ _15169_ _15170_ _14861_ VGND VGND VPWR VPWR _15171_ sky130_fd_sc_hd__a22o_1
X_18413_ registers\[56\]\[1\] registers\[57\]\[1\] registers\[58\]\[1\] registers\[59\]\[1\]
+ _05079_ _05081_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux4_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31671_ _14342_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19393_ registers\[44\]\[29\] registers\[45\]\[29\] registers\[46\]\[29\] registers\[47\]\[29\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux4_1
XFILLER_37_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33410_ clknet_leaf_256_CLK _01524_ VGND VGND VPWR VPWR registers\[46\]\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _05039_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__buf_4
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30622_ _13779_ VGND VGND VPWR VPWR _13791_ sky130_fd_sc_hd__buf_4
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34390_ clknet_leaf_94_CLK _02504_ VGND VGND VPWR VPWR registers\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33341_ clknet_leaf_274_CLK _01455_ VGND VGND VPWR VPWR registers\[47\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_18275_ net79 net80 VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__nor2b_4
XFILLER_175_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30553_ _09778_ registers\[13\]\[41\] _13753_ VGND VGND VPWR VPWR _13755_ sky130_fd_sc_hd__mux2_1
XFILLER_202_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17226_ _14578_ VGND VGND VPWR VPWR _15708_ sky130_fd_sc_hd__buf_4
X_36060_ clknet_leaf_37_CLK _04174_ VGND VGND VPWR VPWR registers\[59\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33272_ clknet_leaf_336_CLK _01386_ VGND VGND VPWR VPWR registers\[48\]\[42\] sky130_fd_sc_hd__dfxtp_1
Xinput10 DW[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_6
XFILLER_175_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30484_ _13718_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__clkbuf_1
Xinput21 DW[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput32 DW[38] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
XFILLER_204_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35011_ clknet_leaf_204_CLK _03125_ VGND VGND VPWR VPWR registers\[21\]\[53\] sky130_fd_sc_hd__dfxtp_1
Xinput43 DW[48] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_6
XFILLER_239_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32223_ clknet_leaf_240_CLK _00337_ VGND VGND VPWR VPWR registers\[9\]\[54\] sky130_fd_sc_hd__dfxtp_1
Xinput54 DW[58] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_12
X_17157_ _14607_ VGND VGND VPWR VPWR _15641_ sky130_fd_sc_hd__buf_4
Xinput65 R1[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput76 R2[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput87 RW[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_239_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16108_ _14571_ VGND VGND VPWR VPWR _14621_ sky130_fd_sc_hd__clkbuf_8
XFILLER_196_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32154_ clknet_leaf_24_CLK _00268_ VGND VGND VPWR VPWR registers\[39\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17088_ registers\[40\]\[29\] registers\[41\]\[29\] registers\[42\]\[29\] registers\[43\]\[29\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15573_ sky130_fd_sc_hd__mux4_1
XFILLER_131_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31105_ registers\[0\]\[47\] _13033_ _14037_ VGND VGND VPWR VPWR _14045_ sky130_fd_sc_hd__mux2_1
XFILLER_83_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16039_ net69 VGND VGND VPWR VPWR _14553_ sky130_fd_sc_hd__buf_12
XFILLER_100_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32085_ clknet_leaf_490_CLK _00061_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_30_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_30_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35913_ clknet_leaf_160_CLK _04027_ VGND VGND VPWR VPWR registers\[7\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_31036_ registers\[0\]\[14\] _12964_ _14004_ VGND VGND VPWR VPWR _14009_ sky130_fd_sc_hd__mux2_1
XFILLER_233_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35844_ clknet_leaf_226_CLK _03958_ VGND VGND VPWR VPWR registers\[8\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_59__f_CLK clknet_5_29_0_CLK VGND VGND VPWR VPWR clknet_6_59__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_211_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19729_ registers\[4\]\[38\] registers\[5\]\[38\] registers\[6\]\[38\] registers\[7\]\[38\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux4_1
X_35775_ clknet_leaf_300_CLK _03889_ VGND VGND VPWR VPWR registers\[0\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_32987_ clknet_leaf_52_CLK _01101_ VGND VGND VPWR VPWR registers\[52\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22740_ registers\[0\]\[59\] registers\[1\]\[59\] registers\[2\]\[59\] registers\[3\]\[59\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__mux4_1
X_34726_ clknet_leaf_451_CLK _02840_ VGND VGND VPWR VPWR registers\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31938_ _09815_ registers\[49\]\[58\] _14474_ VGND VGND VPWR VPWR _14483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22671_ _09309_ _09312_ _09083_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__o21ba_1
XFILLER_168_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34657_ clknet_leaf_9_CLK _02771_ VGND VGND VPWR VPWR registers\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31869_ _09742_ registers\[49\]\[25\] _14441_ VGND VGND VPWR VPWR _14447_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_97_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_97_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24410_ net49 VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__buf_4
XFILLER_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21622_ registers\[36\]\[27\] registers\[37\]\[27\] registers\[38\]\[27\] registers\[39\]\[27\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__mux4_1
XFILLER_94_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33608_ clknet_leaf_243_CLK _01722_ VGND VGND VPWR VPWR registers\[43\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25390_ _10793_ registers\[50\]\[30\] _10970_ VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__mux2_1
XFILLER_21_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34588_ clknet_leaf_4_CLK _02702_ VGND VGND VPWR VPWR registers\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24341_ _10369_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
X_21553_ registers\[56\]\[25\] registers\[57\]\[25\] registers\[58\]\[25\] registers\[59\]\[25\]
+ _08194_ _07984_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__mux4_1
X_33539_ clknet_leaf_255_CLK _01653_ VGND VGND VPWR VPWR registers\[44\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20504_ _05060_ _07204_ _07205_ _05066_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__a22o_1
XFILLER_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24272_ _10322_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27060_ _11767_ registers\[38\]\[18\] _11876_ VGND VGND VPWR VPWR _11885_ sky130_fd_sc_hd__mux2_1
X_21484_ registers\[36\]\[23\] registers\[37\]\[23\] registers\[38\]\[23\] registers\[39\]\[23\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__mux4_1
XFILLER_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26011_ _10728_ registers\[45\]\[0\] _11301_ VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__mux2_1
X_23223_ net19 VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__clkbuf_4
X_35209_ clknet_leaf_155_CLK _03323_ VGND VGND VPWR VPWR registers\[18\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20435_ registers\[60\]\[59\] registers\[61\]\[59\] registers\[62\]\[59\] registers\[63\]\[59\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__mux4_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36189_ clknet_leaf_93_CLK _00070_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_1
XFILLER_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23154_ _09703_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XTAP_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20366_ registers\[32\]\[57\] registers\[33\]\[57\] registers\[34\]\[57\] registers\[35\]\[57\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__mux4_1
XFILLER_173_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22105_ _07352_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__buf_4
XTAP_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23085_ _09655_ VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__buf_6
XTAP_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27962_ registers\[32\]\[61\] _10432_ _12292_ VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__mux2_1
X_20297_ registers\[16\]\[54\] registers\[17\]\[54\] registers\[18\]\[54\] registers\[19\]\[54\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_21_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_21_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29701_ _13306_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__clkbuf_1
XTAP_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26913_ _11790_ registers\[3\]\[29\] _11772_ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__mux2_1
X_22036_ registers\[20\]\[38\] registers\[21\]\[38\] registers\[22\]\[38\] registers\[23\]\[38\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__mux4_1
XTAP_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27893_ registers\[32\]\[28\] _10363_ _12315_ VGND VGND VPWR VPWR _12324_ sky130_fd_sc_hd__mux2_1
XFILLER_248_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29632_ registers\[20\]\[53\] _13046_ _13266_ VGND VGND VPWR VPWR _13270_ sky130_fd_sc_hd__mux2_1
XTAP_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26844_ net62 VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29563_ registers\[20\]\[20\] _12976_ _13233_ VGND VGND VPWR VPWR _13234_ sky130_fd_sc_hd__mux2_1
XFILLER_180_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26775_ _11704_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__clkbuf_1
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23987_ _09527_ registers\[5\]\[6\] _10161_ VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28514_ _11734_ registers\[27\]\[2\] _12648_ VGND VGND VPWR VPWR _12651_ sky130_fd_sc_hd__mux2_1
XFILLER_217_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25726_ _11150_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29494_ _13197_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22938_ net11 VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28445_ _12614_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25657_ _11114_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
X_22869_ registers\[28\]\[63\] registers\[29\]\[63\] registers\[30\]\[63\] registers\[31\]\[63\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__mux4_1
XFILLER_188_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_88_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24608_ _10527_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16390_ _14891_ _14894_ _14525_ VGND VGND VPWR VPWR _14895_ sky130_fd_sc_hd__o21ba_2
X_28376_ _12578_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_1
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25588_ _11076_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27327_ _12025_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__clkbuf_1
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24539_ _10489_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18060_ registers\[20\]\[56\] registers\[21\]\[56\] registers\[22\]\[56\] registers\[23\]\[56\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux4_1
XFILLER_157_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27258_ _11830_ registers\[37\]\[48\] _11980_ VGND VGND VPWR VPWR _11989_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17011_ registers\[20\]\[26\] registers\[21\]\[26\] registers\[22\]\[26\] registers\[23\]\[26\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15499_ sky130_fd_sc_hd__mux4_1
X_26209_ _10793_ registers\[44\]\[30\] _11405_ VGND VGND VPWR VPWR _11406_ sky130_fd_sc_hd__mux2_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27189_ _11761_ registers\[37\]\[15\] _11947_ VGND VGND VPWR VPWR _11953_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18962_ _05708_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_12_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_12_CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_1600 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1611 _15105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17913_ _04682_ _04687_ _04611_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1622 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1633 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18893_ registers\[40\]\[15\] registers\[41\]\[15\] registers\[42\]\[15\] registers\[43\]\[15\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__mux4_1
XTAP_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1644 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1655 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1666 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ _04615_ _04618_ _04619_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__o211a_1
X_32910_ clknet_leaf_179_CLK _01024_ VGND VGND VPWR VPWR registers\[53\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1677 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33890_ clknet_leaf_47_CLK _02004_ VGND VGND VPWR VPWR registers\[38\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1688 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1699 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32841_ clknet_leaf_177_CLK _00955_ VGND VGND VPWR VPWR registers\[55\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17775_ _04547_ _04553_ _15963_ _15964_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__o211a_1
XFILLER_66_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19514_ _06241_ _06244_ _06169_ _06170_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__o211a_1
X_16726_ registers\[24\]\[18\] registers\[25\]\[18\] registers\[26\]\[18\] registers\[27\]\[18\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15222_ sky130_fd_sc_hd__mux4_1
X_32772_ clknet_leaf_234_CLK _00886_ VGND VGND VPWR VPWR registers\[56\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_35560_ clknet_leaf_398_CLK _03674_ VGND VGND VPWR VPWR registers\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34511_ clknet_leaf_111_CLK _02625_ VGND VGND VPWR VPWR registers\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_19445_ registers\[4\]\[30\] registers\[5\]\[30\] registers\[6\]\[30\] registers\[7\]\[30\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__mux4_1
X_31723_ _14347_ VGND VGND VPWR VPWR _14370_ sky130_fd_sc_hd__buf_4
X_16657_ registers\[28\]\[16\] registers\[29\]\[16\] registers\[30\]\[16\] registers\[31\]\[16\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15155_ sky130_fd_sc_hd__mux4_1
X_35491_ clknet_leaf_469_CLK _03605_ VGND VGND VPWR VPWR registers\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_79_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_223_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34442_ clknet_leaf_166_CLK _02556_ VGND VGND VPWR VPWR registers\[30\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_31654_ registers\[63\]\[51\] net47 _14332_ VGND VGND VPWR VPWR _14334_ sky130_fd_sc_hd__mux2_1
X_19376_ registers\[4\]\[28\] registers\[5\]\[28\] registers\[6\]\[28\] registers\[7\]\[28\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__mux4_1
XFILLER_206_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16588_ registers\[20\]\[14\] registers\[21\]\[14\] registers\[22\]\[14\] registers\[23\]\[14\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15088_ sky130_fd_sc_hd__mux4_1
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30605_ _13782_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__clkbuf_1
X_18327_ _05041_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__buf_12
XFILLER_148_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34373_ clknet_leaf_213_CLK _02487_ VGND VGND VPWR VPWR registers\[31\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31585_ _14297_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_945 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36112_ clknet_leaf_75_CLK _04226_ VGND VGND VPWR VPWR registers\[49\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_33324_ clknet_leaf_345_CLK _01438_ VGND VGND VPWR VPWR registers\[47\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_18258_ _05018_ _05021_ _14553_ _14555_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__o211a_1
X_30536_ _09760_ registers\[13\]\[33\] _13742_ VGND VGND VPWR VPWR _13746_ sky130_fd_sc_hd__mux2_1
XFILLER_129_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17209_ registers\[48\]\[32\] registers\[49\]\[32\] registers\[50\]\[32\] registers\[51\]\[32\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15691_ sky130_fd_sc_hd__mux4_1
X_36043_ clknet_leaf_167_CLK _04157_ VGND VGND VPWR VPWR registers\[63\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33255_ clknet_leaf_436_CLK _01369_ VGND VGND VPWR VPWR registers\[48\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30467_ _09648_ registers\[13\]\[0\] _13709_ VGND VGND VPWR VPWR _13710_ sky130_fd_sc_hd__mux2_1
X_18189_ registers\[36\]\[61\] registers\[37\]\[61\] registers\[38\]\[61\] registers\[39\]\[61\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux4_1
XFILLER_116_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20220_ _06927_ _06930_ _06855_ _06856_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__o211a_1
XFILLER_144_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32206_ clknet_leaf_415_CLK _00320_ VGND VGND VPWR VPWR registers\[9\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33186_ clknet_leaf_469_CLK _01300_ VGND VGND VPWR VPWR registers\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_30398_ _13673_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__clkbuf_1
X_20151_ registers\[4\]\[50\] registers\[5\]\[50\] registers\[6\]\[50\] registers\[7\]\[50\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__mux4_1
X_32137_ clknet_leaf_397_CLK _00054_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32068_ clknet_leaf_202_CLK _00246_ VGND VGND VPWR VPWR registers\[62\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_20082_ registers\[4\]\[48\] registers\[5\]\[48\] registers\[6\]\[48\] registers\[7\]\[48\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux4_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31019_ registers\[0\]\[6\] _12947_ _13993_ VGND VGND VPWR VPWR _14000_ sky130_fd_sc_hd__mux2_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _09586_ registers\[60\]\[34\] _10122_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__mux2_1
XFILLER_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24890_ _10676_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23841_ _09517_ registers\[60\]\[1\] _10089_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__mux2_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35827_ clknet_leaf_383_CLK _03941_ VGND VGND VPWR VPWR registers\[8\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26560_ _10739_ registers\[41\]\[4\] _11586_ VGND VGND VPWR VPWR _11591_ sky130_fd_sc_hd__mux2_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_508 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20984_ _07305_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__clkbuf_8
X_35758_ clknet_leaf_377_CLK _03872_ VGND VGND VPWR VPWR registers\[0\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_23772_ _09584_ registers\[29\]\[33\] _10050_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__mux2_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_519 _00168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25511_ _11036_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_1
X_22723_ _09342_ _09349_ _09356_ _09363_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__or4_4
X_34709_ clknet_leaf_95_CLK _02823_ VGND VGND VPWR VPWR registers\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26491_ _10806_ registers\[42\]\[36\] _11547_ VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__mux2_1
X_35689_ clknet_leaf_460_CLK _03803_ VGND VGND VPWR VPWR registers\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_28230_ _11855_ registers\[30\]\[60\] _12434_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__mux2_1
X_25442_ _10846_ registers\[50\]\[55\] _10992_ VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22654_ _07296_ _09295_ _09296_ _07302_ VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__a22o_1
XFILLER_186_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28161_ _11786_ registers\[30\]\[27\] _12457_ VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__mux2_1
X_21605_ registers\[24\]\[26\] registers\[25\]\[26\] registers\[26\]\[26\] registers\[27\]\[26\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__mux4_1
X_22585_ _09020_ _09228_ _09229_ _09024_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__a22o_1
XFILLER_51_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25373_ _10777_ registers\[50\]\[22\] _10959_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__mux2_1
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27112_ _11912_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24324_ registers\[57\]\[25\] _10357_ _10347_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__mux2_1
X_28092_ _12428_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__clkbuf_1
X_21536_ _07349_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__buf_4
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27043_ _11864_ VGND VGND VPWR VPWR _11876_ sky130_fd_sc_hd__buf_6
X_24255_ net34 VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__buf_4
X_21467_ _07929_ _08142_ _08143_ _07932_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__a22o_1
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20418_ _06868_ _07121_ _07122_ _06871_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__a22o_1
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23206_ registers\[9\]\[19\] _09697_ _09722_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__mux2_1
XFILLER_175_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24186_ _09590_ registers\[58\]\[36\] _10266_ VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__mux2_1
X_21398_ registers\[16\]\[20\] registers\[17\]\[20\] registers\[18\]\[20\] registers\[19\]\[20\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__mux4_1
XFILLER_190_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20349_ registers\[8\]\[56\] registers\[9\]\[56\] registers\[10\]\[56\] registers\[11\]\[56\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__mux4_1
X_23137_ registers\[39\]\[16\] _09691_ _09679_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__mux2_1
XTAP_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28994_ registers\[24\]\[38\] _10384_ _12894_ VGND VGND VPWR VPWR _12903_ sky130_fd_sc_hd__mux2_1
XTAP_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27945_ _12351_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__clkbuf_1
X_23068_ net58 VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__buf_2
XTAP_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22019_ registers\[52\]\[38\] registers\[53\]\[38\] registers\[54\]\[38\] registers\[55\]\[38\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__mux4_1
XTAP_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27876_ _12292_ VGND VGND VPWR VPWR _12315_ sky130_fd_sc_hd__buf_4
XFILLER_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26827_ _11732_ registers\[3\]\[1\] _11730_ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__mux2_1
XTAP_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29615_ registers\[20\]\[45\] _13029_ _13255_ VGND VGND VPWR VPWR _13261_ sky130_fd_sc_hd__mux2_1
XTAP_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_6_42__f_CLK clknet_5_21_0_CLK VGND VGND VPWR VPWR clknet_6_42__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_229_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _04339_ _04344_ _15955_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__o21ba_1
X_29546_ registers\[20\]\[12\] _12960_ _13222_ VGND VGND VPWR VPWR _13225_ sky130_fd_sc_hd__mux2_1
XFILLER_75_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26758_ _11695_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16511_ _14796_ _15011_ _15012_ _14799_ VGND VGND VPWR VPWR _15013_ sky130_fd_sc_hd__a22o_1
X_25709_ registers\[48\]\[50\] _10409_ _11141_ VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__mux2_1
X_29477_ _13188_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17491_ _15959_ _15962_ _15963_ _15964_ VGND VGND VPWR VPWR _15965_ sky130_fd_sc_hd__o211a_1
X_26689_ _11659_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_868 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19230_ _05688_ _05967_ _05968_ _05691_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a22o_1
X_28428_ _12605_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__clkbuf_1
X_16442_ _14941_ _14944_ _14945_ VGND VGND VPWR VPWR _14946_ sky130_fd_sc_hd__o21ba_1
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_1_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_220_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19161_ _05898_ _05901_ _05826_ _05827_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__o211a_1
X_28359_ registers\[2\]\[57\] _10424_ _12561_ VGND VGND VPWR VPWR _12569_ sky130_fd_sc_hd__mux2_1
X_16373_ registers\[24\]\[8\] registers\[25\]\[8\] registers\[26\]\[8\] registers\[27\]\[8\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14879_ sky130_fd_sc_hd__mux4_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18112_ registers\[12\]\[58\] registers\[13\]\[58\] registers\[14\]\[58\] registers\[15\]\[58\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__mux4_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31370_ _14184_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__clkbuf_1
X_19092_ registers\[4\]\[20\] registers\[5\]\[20\] registers\[6\]\[20\] registers\[7\]\[20\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__mux4_1
XFILLER_219_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30321_ registers\[15\]\[60\] _13060_ _13565_ VGND VGND VPWR VPWR _13632_ sky130_fd_sc_hd__mux2_1
X_18043_ registers\[48\]\[56\] registers\[49\]\[56\] registers\[50\]\[56\] registers\[51\]\[56\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux4_1
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33040_ clknet_leaf_75_CLK _01154_ VGND VGND VPWR VPWR registers\[51\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_30252_ registers\[15\]\[27\] _12991_ _13588_ VGND VGND VPWR VPWR _13596_ sky130_fd_sc_hd__mux2_1
XFILLER_153_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30183_ _13559_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19994_ registers\[60\]\[46\] registers\[61\]\[46\] registers\[62\]\[46\] registers\[63\]\[46\]
+ _06648_ _06442_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__mux4_1
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18945_ _05688_ _05689_ _05690_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a22o_1
XFILLER_80_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34991_ clknet_leaf_387_CLK _03105_ VGND VGND VPWR VPWR registers\[21\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1430 _05008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1441 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1452 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33942_ clknet_leaf_120_CLK _02056_ VGND VGND VPWR VPWR registers\[37\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1463 _05159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1474 _05466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18876_ registers\[0\]\[14\] registers\[1\]\[14\] registers\[2\]\[14\] registers\[3\]\[14\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__mux4_1
XTAP_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1485 _06807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1496 _07324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17827_ registers\[32\]\[50\] registers\[33\]\[50\] registers\[34\]\[50\] registers\[35\]\[50\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__mux4_1
X_33873_ clknet_leaf_134_CLK _01987_ VGND VGND VPWR VPWR registers\[38\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35612_ clknet_leaf_15_CLK _03726_ VGND VGND VPWR VPWR registers\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_32824_ clknet_leaf_331_CLK _00938_ VGND VGND VPWR VPWR registers\[55\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_17758_ registers\[36\]\[48\] registers\[37\]\[48\] registers\[38\]\[48\] registers\[39\]\[48\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__mux4_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35543_ clknet_leaf_81_CLK _03657_ VGND VGND VPWR VPWR registers\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16709_ _15198_ _15200_ _15203_ _15204_ VGND VGND VPWR VPWR _15205_ sky130_fd_sc_hd__a22o_1
X_17689_ _04340_ _04468_ _04469_ _04343_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a22o_1
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32755_ clknet_leaf_363_CLK _00869_ VGND VGND VPWR VPWR registers\[56\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31706_ _14361_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__clkbuf_1
X_19428_ _05073_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__buf_2
X_35474_ clknet_leaf_77_CLK _03588_ VGND VGND VPWR VPWR registers\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32686_ clknet_leaf_371_CLK _00800_ VGND VGND VPWR VPWR registers\[57\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34425_ clknet_leaf_60_CLK _02539_ VGND VGND VPWR VPWR registers\[30\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31637_ registers\[63\]\[43\] net38 _14321_ VGND VGND VPWR VPWR _14325_ sky130_fd_sc_hd__mux2_1
X_19359_ _05092_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__clkbuf_8
XFILLER_91_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22370_ _07328_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__buf_4
XFILLER_241_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31568_ registers\[63\]\[10\] net2 _14288_ VGND VGND VPWR VPWR _14289_ sky130_fd_sc_hd__mux2_1
X_34356_ clknet_leaf_416_CLK _02470_ VGND VGND VPWR VPWR registers\[31\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21321_ _07361_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__buf_6
XFILLER_191_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33307_ clknet_leaf_31_CLK _01421_ VGND VGND VPWR VPWR registers\[47\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_30519_ _09742_ registers\[13\]\[25\] _13731_ VGND VGND VPWR VPWR _13737_ sky130_fd_sc_hd__mux2_1
X_34287_ clknet_leaf_352_CLK _02401_ VGND VGND VPWR VPWR registers\[32\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31499_ _14252_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33238_ clknet_leaf_69_CLK _01352_ VGND VGND VPWR VPWR registers\[48\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_36026_ clknet_leaf_287_CLK _04140_ VGND VGND VPWR VPWR registers\[63\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_24040_ _09580_ registers\[5\]\[31\] _10194_ VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__mux2_1
X_21252_ registers\[24\]\[16\] registers\[25\]\[16\] registers\[26\]\[16\] registers\[27\]\[16\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__mux4_1
XFILLER_116_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20203_ _05045_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__buf_6
XFILLER_172_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33169_ clknet_leaf_76_CLK _01283_ VGND VGND VPWR VPWR registers\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21183_ _07349_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__buf_4
XFILLER_145_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20134_ _05073_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__buf_2
XFILLER_89_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25991_ _10846_ registers\[46\]\[55\] _11285_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27730_ _12238_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__clkbuf_1
X_20065_ _05092_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__clkbuf_4
X_24942_ _09601_ registers\[53\]\[41\] _10702_ VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__mux2_1
XFILLER_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27661_ registers\[34\]\[46\] _10401_ _12195_ VGND VGND VPWR VPWR _12202_ sky130_fd_sc_hd__mux2_1
XFILLER_86_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24873_ _10667_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29400_ _09672_ registers\[21\]\[7\] _13140_ VGND VGND VPWR VPWR _13148_ sky130_fd_sc_hd__mux2_1
XFILLER_39_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26612_ _10791_ registers\[41\]\[29\] _11608_ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__mux2_1
X_23824_ _09636_ registers\[29\]\[58\] _10072_ VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27592_ registers\[34\]\[13\] _10332_ _12162_ VGND VGND VPWR VPWR _12166_ sky130_fd_sc_hd__mux2_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_327 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29331_ _13111_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26543_ _10858_ registers\[42\]\[61\] _11513_ VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__mux2_1
XFILLER_214_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_338 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23755_ _09567_ registers\[29\]\[25\] _10039_ VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__mux2_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_349 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20967_ registers\[12\]\[8\] registers\[13\]\[8\] registers\[14\]\[8\] registers\[15\]\[8\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__mux4_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22706_ registers\[52\]\[58\] registers\[53\]\[58\] registers\[54\]\[58\] registers\[55\]\[58\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__mux4_1
X_29262_ _13075_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26474_ _10789_ registers\[42\]\[28\] _11536_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__mux2_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23686_ registers\[61\]\[58\] _09815_ _09998_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__mux2_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _07585_ _07590_ _07370_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__o21ba_1
X_28213_ _12492_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25425_ _10829_ registers\[50\]\[47\] _10981_ VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__mux2_1
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22637_ _09148_ _09278_ _09279_ _09153_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__a22o_1
XFILLER_213_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29193_ _13030_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28144_ _11769_ registers\[30\]\[19\] _12446_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__mux2_1
XFILLER_70_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25356_ _10760_ registers\[50\]\[14\] _10948_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__mux2_1
XFILLER_22_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22568_ _09210_ _09213_ _09116_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__o21ba_1
XFILLER_210_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24307_ net13 VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__buf_4
X_28075_ _11834_ registers\[31\]\[50\] _12419_ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__mux2_1
X_21519_ _07314_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__buf_6
XFILLER_182_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25287_ _10827_ registers\[51\]\[46\] _10909_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__mux2_1
X_22499_ _09125_ _09132_ _09139_ _09146_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__or4_4
XFILLER_181_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27026_ _11867_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__clkbuf_1
X_24238_ _09642_ registers\[58\]\[61\] _10232_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__mux2_1
XFILLER_135_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24169_ _09573_ registers\[58\]\[28\] _10255_ VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__mux2_1
XFILLER_150_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16991_ registers\[52\]\[26\] registers\[53\]\[26\] registers\[54\]\[26\] registers\[55\]\[26\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15479_ sky130_fd_sc_hd__mux4_1
XFILLER_205_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28977_ net282 VGND VGND VPWR VPWR _12894_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18730_ _05102_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__buf_4
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27928_ _12342_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _05065_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__buf_4
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27859_ _12306_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__clkbuf_1
XTAP_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ registers\[28\]\[43\] registers\[29\]\[43\] registers\[30\]\[43\] registers\[31\]\[43\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__mux4_1
X_30870_ _09705_ _12149_ VGND VGND VPWR VPWR _13921_ sky130_fd_sc_hd__nor2_8
XFILLER_218_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _05345_ _05346_ _05347_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__a22o_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17543_ registers\[20\]\[41\] registers\[21\]\[41\] registers\[22\]\[41\] registers\[23\]\[41\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__mux4_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29529_ registers\[20\]\[4\] _12943_ _13211_ VGND VGND VPWR VPWR _13216_ sky130_fd_sc_hd__mux2_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_850 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_861 _09306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32540_ clknet_leaf_477_CLK _00654_ VGND VGND VPWR VPWR registers\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_872 _09510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17474_ registers\[32\]\[40\] registers\[33\]\[40\] registers\[34\]\[40\] registers\[35\]\[40\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _15948_ sky130_fd_sc_hd__mux4_1
XFILLER_220_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_883 _09580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_894 _09648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ registers\[48\]\[10\] registers\[49\]\[10\] registers\[50\]\[10\] registers\[51\]\[10\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _14929_ sky130_fd_sc_hd__mux4_1
X_19213_ registers\[32\]\[24\] registers\[33\]\[24\] registers\[34\]\[24\] registers\[35\]\[24\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__mux4_1
X_32471_ clknet_leaf_61_CLK _00585_ VGND VGND VPWR VPWR registers\[60\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31422_ _09668_ registers\[6\]\[5\] _14206_ VGND VGND VPWR VPWR _14212_ sky130_fd_sc_hd__mux2_1
X_34210_ clknet_leaf_56_CLK _02324_ VGND VGND VPWR VPWR registers\[33\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_19144_ _05045_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__buf_4
X_16356_ _14855_ _14857_ _14860_ _14861_ VGND VGND VPWR VPWR _14862_ sky130_fd_sc_hd__a22o_1
X_35190_ clknet_leaf_310_CLK _03304_ VGND VGND VPWR VPWR registers\[18\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34141_ clknet_leaf_22_CLK _02255_ VGND VGND VPWR VPWR registers\[34\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_31353_ _14175_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__clkbuf_1
X_19075_ _05073_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__buf_2
XFILLER_185_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16287_ _14789_ _14794_ _14554_ _14556_ VGND VGND VPWR VPWR _14795_ sky130_fd_sc_hd__o211a_1
XFILLER_199_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18026_ registers\[24\]\[55\] registers\[25\]\[55\] registers\[26\]\[55\] registers\[27\]\[55\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__mux4_1
X_30304_ _13623_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34072_ clknet_leaf_34_CLK _02186_ VGND VGND VPWR VPWR registers\[35\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_31284_ _14139_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33023_ clknet_leaf_268_CLK _01137_ VGND VGND VPWR VPWR registers\[52\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_30235_ registers\[15\]\[19\] _12974_ _13577_ VGND VGND VPWR VPWR _13587_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30166_ registers\[16\]\[50\] _13039_ _13550_ VGND VGND VPWR VPWR _13551_ sky130_fd_sc_hd__mux2_1
XFILLER_114_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19977_ _06525_ _06693_ _06694_ _06528_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__a22o_1
XFILLER_115_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18928_ registers\[44\]\[16\] registers\[45\]\[16\] registers\[46\]\[16\] registers\[47\]\[16\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__mux4_1
X_34974_ clknet_leaf_491_CLK _03088_ VGND VGND VPWR VPWR registers\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30097_ _13514_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1260 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1271 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1282 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33925_ clknet_leaf_261_CLK _02039_ VGND VGND VPWR VPWR registers\[38\]\[55\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1293 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18859_ registers\[40\]\[14\] registers\[41\]\[14\] registers\[42\]\[14\] registers\[43\]\[14\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__mux4_1
XFILLER_227_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33856_ clknet_leaf_225_CLK _01970_ VGND VGND VPWR VPWR registers\[3\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21870_ _08469_ _08533_ _08534_ _08472_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__a22o_1
XFILLER_242_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20821_ _07511_ _07515_ _07339_ _07341_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__o211a_1
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32807_ clknet_leaf_438_CLK _00921_ VGND VGND VPWR VPWR registers\[55\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30999_ registers\[10\]\[61\] _13062_ _13921_ VGND VGND VPWR VPWR _13989_ sky130_fd_sc_hd__mux2_1
X_33787_ clknet_leaf_279_CLK _01901_ VGND VGND VPWR VPWR registers\[40\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23540_ _09929_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
X_35526_ clknet_leaf_215_CLK _03640_ VGND VGND VPWR VPWR registers\[13\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20752_ registers\[60\]\[2\] registers\[61\]\[2\] registers\[62\]\[2\] registers\[63\]\[2\]
+ _07327_ _07329_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__mux4_1
X_32738_ clknet_leaf_443_CLK _00852_ VGND VGND VPWR VPWR registers\[56\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35457_ clknet_leaf_238_CLK _03571_ VGND VGND VPWR VPWR registers\[14\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_20683_ _07284_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__buf_12
X_23471_ _09893_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32669_ clknet_leaf_49_CLK _00783_ VGND VGND VPWR VPWR registers\[57\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25210_ _10875_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__clkbuf_1
X_22422_ _08766_ _09070_ _09071_ _08771_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__a22o_1
X_34408_ clknet_leaf_455_CLK _02522_ VGND VGND VPWR VPWR registers\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_26190_ _10775_ registers\[44\]\[21\] _11394_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__mux2_1
X_35388_ clknet_leaf_306_CLK _03502_ VGND VGND VPWR VPWR registers\[15\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25141_ _10831_ registers\[52\]\[48\] _10815_ VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22353_ _09004_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
X_34339_ clknet_leaf_473_CLK _02453_ VGND VGND VPWR VPWR registers\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_6__f_CLK clknet_5_3_0_CLK VGND VGND VPWR VPWR clknet_6_6__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_21304_ registers\[56\]\[18\] registers\[57\]\[18\] registers\[58\]\[18\] registers\[59\]\[18\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__mux4_1
XFILLER_191_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22284_ registers\[40\]\[46\] registers\[41\]\[46\] registers\[42\]\[46\] registers\[43\]\[46\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__mux4_1
X_25072_ net19 VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__buf_2
XFILLER_164_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28900_ _12853_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__clkbuf_1
X_24023_ _09563_ registers\[5\]\[23\] _10183_ VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__mux2_1
X_36009_ clknet_leaf_451_CLK _04123_ VGND VGND VPWR VPWR registers\[63\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_21235_ registers\[60\]\[16\] registers\[61\]\[16\] registers\[62\]\[16\] registers\[63\]\[16\]
+ _07855_ _07649_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__mux4_1
XFILLER_219_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29880_ _13400_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28831_ _12817_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__clkbuf_1
X_21166_ _07314_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__buf_6
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20117_ registers\[24\]\[49\] registers\[25\]\[49\] registers\[26\]\[49\] registers\[27\]\[49\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux4_1
X_28762_ _11847_ registers\[26\]\[56\] _12774_ VGND VGND VPWR VPWR _12781_ sky130_fd_sc_hd__mux2_1
XFILLER_28_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25974_ _10829_ registers\[46\]\[47\] _11274_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__mux2_1
X_21097_ registers\[44\]\[12\] registers\[45\]\[12\] registers\[46\]\[12\] registers\[47\]\[12\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__mux4_1
XFILLER_63_1374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27713_ _12229_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20048_ registers\[28\]\[47\] registers\[29\]\[47\] registers\[30\]\[47\] registers\[31\]\[47\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__mux4_1
X_24925_ _09584_ registers\[53\]\[33\] _10691_ VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28693_ _11778_ registers\[26\]\[23\] _12741_ VGND VGND VPWR VPWR _12745_ sky130_fd_sc_hd__mux2_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27644_ registers\[34\]\[38\] _10384_ _12184_ VGND VGND VPWR VPWR _12193_ sky130_fd_sc_hd__mux2_1
X_24856_ _09510_ registers\[53\]\[0\] _10658_ VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__mux2_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23807_ _10016_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__buf_4
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27575_ registers\[34\]\[5\] _10315_ _12151_ VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__mux2_1
XANTENNA_124 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24787_ _10622_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21999_ _08639_ _08646_ _08653_ _08660_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__or4_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29314_ _09753_ registers\[22\]\[30\] _13102_ VGND VGND VPWR VPWR _13103_ sky130_fd_sc_hd__mux2_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26526_ _11572_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23738_ _09550_ registers\[29\]\[17\] _10028_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__mux2_1
XANTENNA_168 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_179 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29245_ _13065_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__clkbuf_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26457_ _11513_ VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23669_ _09942_ VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__clkbuf_8
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16210_ registers\[36\]\[4\] registers\[37\]\[4\] registers\[38\]\[4\] registers\[39\]\[4\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14720_ sky130_fd_sc_hd__mux4_1
X_25408_ _10812_ registers\[50\]\[39\] _10970_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__mux2_1
X_29176_ _12934_ VGND VGND VPWR VPWR _13019_ sky130_fd_sc_hd__buf_4
X_17190_ registers\[20\]\[31\] registers\[21\]\[31\] registers\[22\]\[31\] registers\[23\]\[31\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15673_ sky130_fd_sc_hd__mux4_1
X_26388_ _10838_ registers\[43\]\[51\] _11498_ VGND VGND VPWR VPWR _11500_ sky130_fd_sc_hd__mux2_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16141_ _14567_ VGND VGND VPWR VPWR _14653_ sky130_fd_sc_hd__buf_4
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28127_ _12447_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__clkbuf_1
X_25339_ _10743_ registers\[50\]\[6\] _10937_ VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__mux2_1
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16072_ _14569_ _14583_ _14585_ VGND VGND VPWR VPWR _14586_ sky130_fd_sc_hd__o21ba_1
X_28058_ _11818_ registers\[31\]\[42\] _12408_ VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__mux2_1
XFILLER_136_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27009_ _11855_ registers\[3\]\[60\] _11729_ VGND VGND VPWR VPWR _11856_ sky130_fd_sc_hd__mux2_1
X_19900_ registers\[8\]\[43\] registers\[9\]\[43\] registers\[10\]\[43\] registers\[11\]\[43\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__mux4_1
XFILLER_170_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30020_ registers\[17\]\[45\] _13029_ _13468_ VGND VGND VPWR VPWR _13474_ sky130_fd_sc_hd__mux2_1
XFILLER_151_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19831_ _06549_ _06552_ _06512_ _06513_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__o211a_1
XFILLER_116_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19762_ _06379_ _06484_ _06485_ _06382_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__a22o_1
X_16974_ _15295_ _15461_ _15462_ _15300_ VGND VGND VPWR VPWR _15463_ sky130_fd_sc_hd__a22o_1
XFILLER_42_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18713_ _05466_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31971_ clknet_leaf_5_CLK _00141_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
X_19693_ registers\[16\]\[37\] registers\[17\]\[37\] registers\[18\]\[37\] registers\[19\]\[37\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__mux4_1
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 DW[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_6
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_292_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_292_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33710_ clknet_leaf_348_CLK _01824_ VGND VGND VPWR VPWR registers\[41\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_18644_ _05197_ _05397_ _05398_ _05202_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__a22o_1
X_30922_ registers\[10\]\[24\] _12985_ _13944_ VGND VGND VPWR VPWR _13949_ sky130_fd_sc_hd__mux2_1
X_34690_ clknet_leaf_223_CLK _02804_ VGND VGND VPWR VPWR registers\[26\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30853_ _13912_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__clkbuf_1
X_33641_ clknet_leaf_430_CLK _01755_ VGND VGND VPWR VPWR registers\[42\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_18575_ registers\[44\]\[6\] registers\[45\]\[6\] registers\[46\]\[6\] registers\[47\]\[6\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__mux4_1
XFILLER_224_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17526_ registers\[48\]\[41\] registers\[49\]\[41\] registers\[50\]\[41\] registers\[51\]\[41\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__mux4_1
XFILLER_229_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33572_ clknet_leaf_57_CLK _01686_ VGND VGND VPWR VPWR registers\[43\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_30784_ _13876_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_680 _05983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35311_ clknet_leaf_394_CLK _03425_ VGND VGND VPWR VPWR registers\[16\]\[33\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_691 _06807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32523_ clknet_leaf_164_CLK _00637_ VGND VGND VPWR VPWR registers\[60\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17457_ registers\[8\]\[39\] registers\[9\]\[39\] registers\[10\]\[39\] registers\[11\]\[39\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15932_ sky130_fd_sc_hd__mux4_1
XFILLER_75_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16408_ registers\[28\]\[9\] registers\[29\]\[9\] registers\[30\]\[9\] registers\[31\]\[9\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14913_ sky130_fd_sc_hd__mux4_1
X_35242_ clknet_leaf_406_CLK _03356_ VGND VGND VPWR VPWR registers\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_32454_ clknet_leaf_213_CLK _00568_ VGND VGND VPWR VPWR registers\[29\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17388_ registers\[12\]\[37\] registers\[13\]\[37\] registers\[14\]\[37\] registers\[15\]\[37\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _15865_ sky130_fd_sc_hd__mux4_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31405_ _14202_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__clkbuf_1
X_16339_ _14842_ _14845_ _14614_ VGND VGND VPWR VPWR _14846_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19127_ registers\[0\]\[21\] registers\[1\]\[21\] registers\[2\]\[21\] registers\[3\]\[21\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__mux4_1
X_32385_ clknet_leaf_233_CLK _00499_ VGND VGND VPWR VPWR registers\[61\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_35173_ clknet_leaf_446_CLK _03287_ VGND VGND VPWR VPWR registers\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34124_ clknet_leaf_169_CLK _02238_ VGND VGND VPWR VPWR registers\[35\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31336_ _14166_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__clkbuf_1
X_19058_ registers\[24\]\[19\] registers\[25\]\[19\] registers\[26\]\[19\] registers\[27\]\[19\]
+ _05631_ _05632_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__mux4_1
XFILLER_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ registers\[36\]\[55\] registers\[37\]\[55\] registers\[38\]\[55\] registers\[39\]\[55\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux4_1
X_31267_ registers\[8\]\[60\] net57 _14063_ VGND VGND VPWR VPWR _14130_ sky130_fd_sc_hd__mux2_1
X_34055_ clknet_leaf_237_CLK _02169_ VGND VGND VPWR VPWR registers\[36\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21020_ registers\[36\]\[10\] registers\[37\]\[10\] registers\[38\]\[10\] registers\[39\]\[10\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__mux4_1
XFILLER_236_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33006_ clknet_leaf_368_CLK _01120_ VGND VGND VPWR VPWR registers\[52\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_30218_ _13578_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__clkbuf_1
X_31198_ registers\[8\]\[27\] net20 _14086_ VGND VGND VPWR VPWR _14094_ sky130_fd_sc_hd__mux2_1
XFILLER_248_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30149_ registers\[16\]\[42\] _13023_ _13539_ VGND VGND VPWR VPWR _13542_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34957_ clknet_leaf_137_CLK _03071_ VGND VGND VPWR VPWR registers\[22\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_22971_ _09576_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1090 _14518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_283_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_283_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24710_ _10580_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21922_ registers\[24\]\[35\] registers\[25\]\[35\] registers\[26\]\[35\] registers\[27\]\[35\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__mux4_1
X_33908_ clknet_leaf_350_CLK _02022_ VGND VGND VPWR VPWR registers\[38\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25690_ registers\[48\]\[41\] _10391_ _11130_ VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__mux2_1
X_34888_ clknet_leaf_210_CLK _03002_ VGND VGND VPWR VPWR registers\[23\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24641_ _10544_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33839_ clknet_leaf_377_CLK _01953_ VGND VGND VPWR VPWR registers\[3\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_21853_ registers\[4\]\[33\] registers\[5\]\[33\] registers\[6\]\[33\] registers\[7\]\[33\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__mux4_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ _07476_ _07483_ _07492_ _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__or4_2
X_27360_ registers\[36\]\[32\] _10372_ _12040_ VGND VGND VPWR VPWR _12043_ sky130_fd_sc_hd__mux2_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24572_ _10506_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21784_ _08272_ _08450_ _08451_ _08275_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__a22o_1
X_26311_ _11459_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
X_23523_ _09920_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__clkbuf_1
X_35509_ clknet_leaf_323_CLK _03623_ VGND VGND VPWR VPWR registers\[13\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_27291_ _09653_ _11010_ VGND VGND VPWR VPWR _12006_ sky130_fd_sc_hd__nor2_8
X_20735_ _07432_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29030_ registers\[24\]\[55\] _10420_ _12916_ VGND VGND VPWR VPWR _12922_ sky130_fd_sc_hd__mux2_1
XFILLER_211_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26242_ _10827_ registers\[44\]\[46\] _11416_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__mux2_1
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23454_ _09884_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20666_ registers\[4\]\[0\] registers\[5\]\[0\] registers\[6\]\[0\] registers\[7\]\[0\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__mux4_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22405_ _09012_ _09053_ _09054_ _09018_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__a22o_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26173_ _10758_ registers\[44\]\[13\] _11383_ VGND VGND VPWR VPWR _11387_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20597_ _07295_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__buf_4
XFILLER_178_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23385_ _09846_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25124_ _10820_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__clkbuf_1
X_22336_ _08677_ _08986_ _08987_ _08681_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__a22o_1
XFILLER_30_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29932_ registers\[17\]\[3\] _12941_ _13424_ VGND VGND VPWR VPWR _13428_ sky130_fd_sc_hd__mux2_1
XFILLER_139_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25055_ _10772_ registers\[52\]\[20\] _10773_ VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__mux2_1
X_22267_ _07289_ VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__buf_4
X_24006_ _09546_ registers\[5\]\[15\] _10172_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__mux2_1
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21218_ _07732_ _07900_ _07901_ _07735_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__a22o_1
X_22198_ _08677_ _08852_ _08853_ _08681_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__a22o_1
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29863_ _13391_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28814_ _12808_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__clkbuf_1
X_21149_ _07829_ _07834_ _07730_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__o21ba_1
X_29794_ _13355_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_238_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28745_ _11830_ registers\[26\]\[48\] _12763_ VGND VGND VPWR VPWR _12772_ sky130_fd_sc_hd__mux2_1
X_25957_ _10812_ registers\[46\]\[39\] _11263_ VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_274_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_274_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24908_ _09567_ registers\[53\]\[25\] _10680_ VGND VGND VPWR VPWR _10686_ sky130_fd_sc_hd__mux2_1
X_16690_ registers\[20\]\[17\] registers\[21\]\[17\] registers\[22\]\[17\] registers\[23\]\[17\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15187_ sky130_fd_sc_hd__mux4_1
X_28676_ _11761_ registers\[26\]\[15\] _12730_ VGND VGND VPWR VPWR _12736_ sky130_fd_sc_hd__mux2_1
X_25888_ _10743_ registers\[46\]\[6\] _11230_ VGND VGND VPWR VPWR _11237_ sky130_fd_sc_hd__mux2_1
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_30_0_CLK clknet_2_3_0_CLK VGND VGND VPWR VPWR clknet_5_30_0_CLK sky130_fd_sc_hd__clkbuf_8
X_24839_ _10649_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27627_ _12150_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__buf_4
XFILLER_98_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__buf_6
XFILLER_215_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27558_ _12146_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__clkbuf_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _15549_ _15788_ _15789_ _15553_ VGND VGND VPWR VPWR _15790_ sky130_fd_sc_hd__a22o_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26509_ _11563_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__buf_4
XFILLER_226_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27489_ _12110_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17242_ _15541_ _15721_ _15722_ _15547_ VGND VGND VPWR VPWR _15723_ sky130_fd_sc_hd__a22o_1
X_29228_ net53 VGND VGND VPWR VPWR _13054_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17173_ registers\[48\]\[31\] registers\[49\]\[31\] registers\[50\]\[31\] registers\[51\]\[31\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15656_ sky130_fd_sc_hd__mux4_1
X_29159_ _13007_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16124_ registers\[4\]\[1\] registers\[5\]\[1\] registers\[6\]\[1\] registers\[7\]\[1\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14637_ sky130_fd_sc_hd__mux4_1
X_32170_ clknet_leaf_81_CLK _00284_ VGND VGND VPWR VPWR registers\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31121_ _14053_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__clkbuf_1
X_16055_ _14558_ _14561_ _14566_ _14568_ VGND VGND VPWR VPWR _14569_ sky130_fd_sc_hd__a22o_1
XFILLER_157_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31052_ _14017_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30003_ registers\[17\]\[37\] _13012_ _13457_ VGND VGND VPWR VPWR _13465_ sky130_fd_sc_hd__mux2_1
XFILLER_69_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19814_ _05162_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35860_ clknet_leaf_82_CLK _03974_ VGND VGND VPWR VPWR registers\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34811_ clknet_leaf_304_CLK _02925_ VGND VGND VPWR VPWR registers\[24\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_19745_ _06226_ _06465_ _06468_ _06231_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__a22o_1
X_35791_ clknet_leaf_137_CLK _03905_ VGND VGND VPWR VPWR registers\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16957_ registers\[52\]\[25\] registers\[53\]\[25\] registers\[54\]\[25\] registers\[55\]\[25\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15446_ sky130_fd_sc_hd__mux4_1
XFILLER_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_265_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_265_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34742_ clknet_leaf_312_CLK _02856_ VGND VGND VPWR VPWR registers\[25\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_31954_ clknet_leaf_0_CLK _00172_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
X_19676_ _06233_ _06398_ _06401_ _06236_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__a22o_1
X_16888_ registers\[48\]\[23\] registers\[49\]\[23\] registers\[50\]\[23\] registers\[51\]\[23\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15379_ sky130_fd_sc_hd__mux4_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18627_ registers\[0\]\[7\] registers\[1\]\[7\] registers\[2\]\[7\] registers\[3\]\[7\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__mux4_1
X_30905_ registers\[10\]\[16\] _12968_ _13933_ VGND VGND VPWR VPWR _13940_ sky130_fd_sc_hd__mux2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34673_ clknet_leaf_409_CLK _02787_ VGND VGND VPWR VPWR registers\[26\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31885_ _14455_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33624_ clknet_leaf_90_CLK _01738_ VGND VGND VPWR VPWR registers\[42\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18558_ _05107_ _05314_ _05315_ _05117_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a22o_1
X_30836_ _13903_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17509_ _14530_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__buf_4
XFILLER_33_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33555_ clknet_leaf_127_CLK _01669_ VGND VGND VPWR VPWR registers\[43\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18489_ registers\[0\]\[3\] registers\[1\]\[3\] registers\[2\]\[3\] registers\[3\]\[3\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__mux4_1
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30767_ _13867_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _05089_ _07219_ _07220_ _05100_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__a22o_1
X_32506_ clknet_leaf_287_CLK _00620_ VGND VGND VPWR VPWR registers\[60\]\[44\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_24 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33486_ clknet_leaf_131_CLK _01600_ VGND VGND VPWR VPWR registers\[44\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30698_ registers\[12\]\[46\] _13031_ _13824_ VGND VGND VPWR VPWR _13831_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_46 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_57 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20451_ _06873_ _07153_ _07154_ _06878_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__a22o_1
X_35225_ clknet_leaf_6_CLK _03339_ VGND VGND VPWR VPWR registers\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_68 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_6_19__f_CLK clknet_5_9_0_CLK VGND VGND VPWR VPWR clknet_6_19__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32437_ clknet_leaf_415_CLK _00551_ VGND VGND VPWR VPWR registers\[29\]\[39\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_79 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1086 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20382_ registers\[12\]\[57\] registers\[13\]\[57\] registers\[14\]\[57\] registers\[15\]\[57\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__mux4_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23170_ _09714_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
X_35156_ clknet_leaf_93_CLK _03270_ VGND VGND VPWR VPWR registers\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32368_ clknet_leaf_369_CLK _00482_ VGND VGND VPWR VPWR registers\[61\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34107_ clknet_leaf_281_CLK _02221_ VGND VGND VPWR VPWR registers\[35\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_22121_ registers\[44\]\[41\] registers\[45\]\[41\] registers\[46\]\[41\] registers\[47\]\[41\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__mux4_1
X_31319_ registers\[7\]\[20\] net13 _14157_ VGND VGND VPWR VPWR _14158_ sky130_fd_sc_hd__mux2_1
X_35087_ clknet_leaf_136_CLK _03201_ VGND VGND VPWR VPWR registers\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_32299_ clknet_leaf_408_CLK _00413_ VGND VGND VPWR VPWR registers\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xoutput120 net120 VGND VGND VPWR VPWR D1[37] sky130_fd_sc_hd__buf_2
Xoutput131 net131 VGND VGND VPWR VPWR D1[47] sky130_fd_sc_hd__buf_2
Xoutput142 net142 VGND VGND VPWR VPWR D1[57] sky130_fd_sc_hd__buf_2
XTAP_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22052_ _08669_ _08710_ _08711_ _08675_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__a22o_1
XTAP_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34038_ clknet_leaf_340_CLK _02152_ VGND VGND VPWR VPWR registers\[36\]\[40\] sky130_fd_sc_hd__dfxtp_1
Xoutput153 net153 VGND VGND VPWR VPWR D1[9] sky130_fd_sc_hd__buf_2
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput164 net164 VGND VGND VPWR VPWR D2[19] sky130_fd_sc_hd__buf_2
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput175 net175 VGND VGND VPWR VPWR D2[29] sky130_fd_sc_hd__buf_2
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput186 net186 VGND VGND VPWR VPWR D2[39] sky130_fd_sc_hd__buf_2
Xoutput197 net197 VGND VGND VPWR VPWR D2[49] sky130_fd_sc_hd__buf_2
XTAP_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _07586_ _07691_ _07692_ _07589_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__a22o_1
XTAP_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26860_ net4 VGND VGND VPWR VPWR _11755_ sky130_fd_sc_hd__clkbuf_4
XTAP_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25811_ _11196_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
X_26791_ _11712_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35989_ clknet_leaf_182_CLK _04103_ VGND VGND VPWR VPWR registers\[63\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_256_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_256_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28530_ _12647_ VGND VGND VPWR VPWR _12659_ sky130_fd_sc_hd__buf_4
XFILLER_244_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25742_ _11160_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22954_ net17 VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__buf_2
XFILLER_228_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21905_ _08565_ _08568_ _08397_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__o21ba_1
X_28461_ _11816_ registers\[28\]\[41\] _12621_ VGND VGND VPWR VPWR _12623_ sky130_fd_sc_hd__mux2_1
X_25673_ registers\[48\]\[33\] _10374_ _11119_ VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__mux2_1
X_22885_ _09518_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27412_ registers\[36\]\[57\] _10424_ _12062_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__mux2_1
X_24624_ _10535_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
X_28392_ _12586_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__clkbuf_1
X_21836_ registers\[44\]\[33\] registers\[45\]\[33\] registers\[46\]\[33\] registers\[47\]\[33\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__mux4_1
XFILLER_243_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27343_ registers\[36\]\[24\] _10355_ _12029_ VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__mux2_1
X_24555_ _09624_ registers\[56\]\[52\] _10495_ VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21767_ _08119_ _08433_ _08434_ _08124_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__a22o_1
XFILLER_180_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23506_ _09911_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
X_27274_ _11997_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__clkbuf_1
X_20718_ _07325_ _07414_ _07415_ _07336_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__a22o_1
XFILLER_145_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24486_ _10461_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
X_21698_ registers\[48\]\[29\] registers\[49\]\[29\] registers\[50\]\[29\] registers\[51\]\[29\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__mux4_1
XFILLER_106_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29013_ registers\[24\]\[47\] _10403_ _12905_ VGND VGND VPWR VPWR _12913_ sky130_fd_sc_hd__mux2_1
XFILLER_200_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26225_ _10810_ registers\[44\]\[38\] _11405_ VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__mux2_1
X_23437_ _09875_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20649_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__buf_6
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26156_ _10741_ registers\[44\]\[5\] _11372_ VGND VGND VPWR VPWR _11378_ sky130_fd_sc_hd__mux2_1
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23368_ _09837_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25107_ _10808_ registers\[52\]\[37\] _10794_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__mux2_1
X_22319_ _08968_ _08971_ _08773_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__o21ba_1
X_26087_ _11341_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
X_23299_ _09794_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29915_ _13418_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25038_ net7 VGND VGND VPWR VPWR _10762_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17860_ _14510_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__clkbuf_4
X_29846_ _13382_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16811_ _15304_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
X_29777_ registers\[1\]\[58\] _13056_ _13337_ VGND VGND VPWR VPWR _13346_ sky130_fd_sc_hd__mux2_1
X_17791_ _04566_ _04569_ _04301_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__o21ba_1
XFILLER_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26989_ _11842_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_247_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_247_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19530_ _06255_ _06260_ _06194_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__o21ba_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28728_ _12718_ VGND VGND VPWR VPWR _12763_ sky130_fd_sc_hd__buf_4
X_16742_ _14998_ _15235_ _15236_ _15001_ VGND VGND VPWR VPWR _15237_ sky130_fd_sc_hd__a22o_1
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16673_ registers\[48\]\[17\] registers\[49\]\[17\] registers\[50\]\[17\] registers\[51\]\[17\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15170_ sky130_fd_sc_hd__mux4_1
X_19461_ _05162_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__buf_2
X_28659_ _11744_ registers\[26\]\[7\] _12719_ VGND VGND VPWR VPWR _12727_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1034 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18412_ _05168_ _05173_ _05074_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31670_ registers\[63\]\[59\] net55 _14332_ VGND VGND VPWR VPWR _14342_ sky130_fd_sc_hd__mux2_1
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _05883_ _06122_ _06125_ _05888_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18343_ _05087_ _05101_ _05103_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__o211a_1
X_30621_ _13790_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__clkbuf_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33340_ clknet_leaf_277_CLK _01454_ VGND VGND VPWR VPWR registers\[47\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_18274_ _05037_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30552_ _13754_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17225_ _14576_ VGND VGND VPWR VPWR _15707_ sky130_fd_sc_hd__buf_6
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30483_ _09674_ registers\[13\]\[8\] _13709_ VGND VGND VPWR VPWR _13718_ sky130_fd_sc_hd__mux2_1
Xinput11 DW[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_6
X_33271_ clknet_leaf_335_CLK _01385_ VGND VGND VPWR VPWR registers\[48\]\[41\] sky130_fd_sc_hd__dfxtp_1
Xinput22 DW[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_4
X_35010_ clknet_leaf_204_CLK _03124_ VGND VGND VPWR VPWR registers\[21\]\[52\] sky130_fd_sc_hd__dfxtp_1
Xinput33 DW[39] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_4
X_32222_ clknet_leaf_242_CLK _00336_ VGND VGND VPWR VPWR registers\[9\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput44 DW[49] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_6
X_17156_ _14530_ VGND VGND VPWR VPWR _15640_ sky130_fd_sc_hd__buf_4
XFILLER_196_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput55 DW[59] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_12
Xinput66 R1[1] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput77 R3[0] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16107_ registers\[44\]\[1\] registers\[45\]\[1\] registers\[46\]\[1\] registers\[47\]\[1\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14620_ sky130_fd_sc_hd__mux4_1
XFILLER_143_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput88 RW[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
X_32153_ clknet_leaf_29_CLK _00267_ VGND VGND VPWR VPWR registers\[39\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17087_ _15572_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31104_ _14044_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__clkbuf_1
X_16038_ _14540_ _14545_ _14550_ _14551_ VGND VGND VPWR VPWR _14552_ sky130_fd_sc_hd__a22o_1
X_32084_ clknet_leaf_490_CLK _00060_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_486_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_486_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_237_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35912_ clknet_leaf_160_CLK _04026_ VGND VGND VPWR VPWR registers\[7\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31035_ _14008_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35843_ clknet_leaf_242_CLK _03957_ VGND VGND VPWR VPWR registers\[8\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17989_ _04481_ _04760_ _04761_ _04484_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_123_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_238_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_238_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19728_ _05127_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__buf_4
XFILLER_226_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35774_ clknet_leaf_300_CLK _03888_ VGND VGND VPWR VPWR registers\[0\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_32986_ clknet_leaf_67_CLK _01100_ VGND VGND VPWR VPWR registers\[52\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34725_ clknet_leaf_445_CLK _02839_ VGND VGND VPWR VPWR registers\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_31937_ _14482_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__clkbuf_1
X_19659_ _05141_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__buf_6
XFILLER_93_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22670_ _09155_ _09310_ _09311_ _09158_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34656_ clknet_leaf_3_CLK _02770_ VGND VGND VPWR VPWR registers\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31868_ _14446_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33607_ clknet_leaf_243_CLK _01721_ VGND VGND VPWR VPWR registers\[43\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_21621_ _07358_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__clkbuf_8
X_30819_ _13894_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34587_ clknet_leaf_22_CLK _02701_ VGND VGND VPWR VPWR registers\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_31799_ registers\[59\]\[56\] net52 _14403_ VGND VGND VPWR VPWR _14410_ sky130_fd_sc_hd__mux2_1
XFILLER_179_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_410_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_410_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24340_ registers\[57\]\[30\] _10367_ _10368_ VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__mux2_1
X_33538_ clknet_leaf_256_CLK _01652_ VGND VGND VPWR VPWR registers\[44\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_21552_ _08222_ _08225_ _08054_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__o21ba_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20503_ registers\[4\]\[61\] registers\[5\]\[61\] registers\[6\]\[61\] registers\[7\]\[61\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__mux4_1
XFILLER_193_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24271_ registers\[57\]\[8\] _10321_ _10305_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__mux2_1
X_33469_ clknet_leaf_274_CLK _01583_ VGND VGND VPWR VPWR registers\[45\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_21483_ registers\[44\]\[23\] registers\[45\]\[23\] registers\[46\]\[23\] registers\[47\]\[23\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__mux4_1
XFILLER_140_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26010_ _11300_ VGND VGND VPWR VPWR _11301_ sky130_fd_sc_hd__buf_4
XFILLER_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35208_ clknet_leaf_153_CLK _03322_ VGND VGND VPWR VPWR registers\[18\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23222_ _09743_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
X_20434_ _05136_ _07136_ _07137_ _05146_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__a22o_1
XFILLER_165_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36188_ clknet_leaf_94_CLK _00069_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35139_ clknet_leaf_241_CLK _03253_ VGND VGND VPWR VPWR registers\[1\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_23153_ registers\[39\]\[21\] _09702_ _09700_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365_ registers\[40\]\[57\] registers\[41\]\[57\] registers\[42\]\[57\] registers\[43\]\[57\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__mux4_1
XFILLER_179_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22104_ registers\[16\]\[40\] registers\[17\]\[40\] registers\[18\]\[40\] registers\[19\]\[40\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__mux4_1
XTAP_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20296_ registers\[24\]\[54\] registers\[25\]\[54\] registers\[26\]\[54\] registers\[27\]\[54\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__mux4_1
X_23084_ _09511_ _09654_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__or2_1
X_27961_ _12359_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__clkbuf_1
XTAP_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29700_ registers\[1\]\[21\] _12979_ _13304_ VGND VGND VPWR VPWR _13306_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_477_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_477_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22035_ registers\[28\]\[38\] registers\[29\]\[38\] registers\[30\]\[38\] registers\[31\]\[38\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__mux4_1
X_26912_ net22 VGND VGND VPWR VPWR _11790_ sky130_fd_sc_hd__clkbuf_4
XTAP_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27892_ _12323_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29631_ _13269_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__clkbuf_1
XTAP_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26843_ _11743_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_229_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_229_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29562_ _13210_ VGND VGND VPWR VPWR _13233_ sky130_fd_sc_hd__buf_4
XFILLER_75_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26774_ registers\[40\]\[41\] _10391_ _11702_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__mux2_1
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23986_ _10167_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28513_ _12650_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__clkbuf_1
X_25725_ registers\[48\]\[58\] _10426_ _11141_ VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__mux2_1
XFILLER_17_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22937_ _09553_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29493_ _09800_ registers\[21\]\[51\] _13195_ VGND VGND VPWR VPWR _13197_ sky130_fd_sc_hd__mux2_1
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28444_ _11799_ registers\[28\]\[33\] _12610_ VGND VGND VPWR VPWR _12614_ sky130_fd_sc_hd__mux2_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25656_ registers\[48\]\[25\] _10357_ _11108_ VGND VGND VPWR VPWR _11114_ sky130_fd_sc_hd__mux2_1
X_22868_ _07343_ _09502_ _09503_ _07353_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__a22o_1
XFILLER_231_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24607_ _09538_ registers\[55\]\[11\] _10525_ VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__mux2_1
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28375_ _11728_ registers\[28\]\[0\] _12577_ VGND VGND VPWR VPWR _12578_ sky130_fd_sc_hd__mux2_1
X_21819_ registers\[4\]\[32\] registers\[5\]\[32\] registers\[6\]\[32\] registers\[7\]\[32\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__mux4_1
X_25587_ registers\[4\]\[58\] _10426_ _11067_ VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__mux2_1
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22799_ registers\[8\]\[61\] registers\[9\]\[61\] registers\[10\]\[61\] registers\[11\]\[61\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__mux4_1
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_401_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_401_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27326_ registers\[36\]\[16\] _10338_ _12018_ VGND VGND VPWR VPWR _12025_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1013 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24538_ _09607_ registers\[56\]\[44\] _10484_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27257_ _11988_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__clkbuf_1
X_24469_ _09538_ registers\[56\]\[11\] _10451_ VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17010_ registers\[28\]\[26\] registers\[29\]\[26\] registers\[30\]\[26\] registers\[31\]\[26\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15498_ sky130_fd_sc_hd__mux4_1
X_26208_ _11371_ VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__buf_4
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27188_ _11952_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_810 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26139_ _11368_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18961_ _05678_ _05687_ _05698_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__or4_1
XFILLER_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1601 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_468_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_468_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17912_ _04683_ _04684_ _04685_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__a22o_1
XANTENNA_1612 _15114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1623 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18892_ _05640_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1634 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1645 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1656 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1667 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17843_ _14555_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__clkbuf_4
X_29829_ _13373_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1678 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1689 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32840_ clknet_leaf_178_CLK _00954_ VGND VGND VPWR VPWR registers\[55\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_17774_ _04548_ _04550_ _04551_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a22o_1
XFILLER_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19513_ _06098_ _06242_ _06243_ _06102_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a22o_1
X_16725_ _15215_ _15220_ _14945_ VGND VGND VPWR VPWR _15221_ sky130_fd_sc_hd__o21ba_1
XFILLER_75_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32771_ clknet_leaf_267_CLK _00885_ VGND VGND VPWR VPWR registers\[56\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34510_ clknet_leaf_109_CLK _02624_ VGND VGND VPWR VPWR registers\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_19444_ registers\[12\]\[30\] registers\[13\]\[30\] registers\[14\]\[30\] registers\[15\]\[30\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__mux4_1
X_31722_ _14369_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__clkbuf_1
X_35490_ clknet_leaf_467_CLK _03604_ VGND VGND VPWR VPWR registers\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_16656_ _14947_ _15150_ _15153_ _14950_ VGND VGND VPWR VPWR _15154_ sky130_fd_sc_hd__a22o_1
XFILLER_90_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34441_ clknet_leaf_214_CLK _02555_ VGND VGND VPWR VPWR registers\[30\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31653_ _14333_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__clkbuf_1
X_19375_ _05127_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__buf_4
XFILLER_76_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16587_ registers\[28\]\[14\] registers\[29\]\[14\] registers\[30\]\[14\] registers\[31\]\[14\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15087_ sky130_fd_sc_hd__mux4_1
XFILLER_15_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30604_ registers\[12\]\[1\] _12937_ _13780_ VGND VGND VPWR VPWR _13782_ sky130_fd_sc_hd__mux2_1
X_18326_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__clkbuf_4
X_34372_ clknet_leaf_205_CLK _02486_ VGND VGND VPWR VPWR registers\[31\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31584_ registers\[63\]\[18\] net10 _14288_ VGND VGND VPWR VPWR _14297_ sky130_fd_sc_hd__mux2_1
XFILLER_148_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36111_ clknet_leaf_171_CLK _04225_ VGND VGND VPWR VPWR registers\[49\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1029 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_957 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33323_ clknet_leaf_429_CLK _01437_ VGND VGND VPWR VPWR registers\[47\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_18257_ _14600_ _05019_ _05020_ _14610_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__a22o_1
X_30535_ _13745_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36042_ clknet_leaf_178_CLK _04156_ VGND VGND VPWR VPWR registers\[63\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_17208_ registers\[56\]\[32\] registers\[57\]\[32\] registers\[58\]\[32\] registers\[59\]\[32\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15690_ sky130_fd_sc_hd__mux4_1
X_30466_ _13708_ VGND VGND VPWR VPWR _13709_ sky130_fd_sc_hd__buf_4
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33254_ clknet_leaf_434_CLK _01368_ VGND VGND VPWR VPWR registers\[48\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18188_ registers\[44\]\[61\] registers\[45\]\[61\] registers\[46\]\[61\] registers\[47\]\[61\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux4_1
XFILLER_141_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32205_ clknet_leaf_354_CLK _00319_ VGND VGND VPWR VPWR registers\[9\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17139_ registers\[8\]\[30\] registers\[9\]\[30\] registers\[10\]\[30\] registers\[11\]\[30\]
+ _15449_ _15450_ VGND VGND VPWR VPWR _15623_ sky130_fd_sc_hd__mux4_1
X_33185_ clknet_leaf_470_CLK _01299_ VGND VGND VPWR VPWR registers\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_30397_ _09756_ registers\[14\]\[31\] _13671_ VGND VGND VPWR VPWR _13673_ sky130_fd_sc_hd__mux2_1
X_20150_ registers\[12\]\[50\] registers\[13\]\[50\] registers\[14\]\[50\] registers\[15\]\[50\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__mux4_1
XFILLER_171_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32136_ clknet_leaf_460_CLK _00053_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_459_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_459_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20081_ _05127_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__buf_4
X_32067_ clknet_leaf_294_CLK _00245_ VGND VGND VPWR VPWR registers\[62\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31018_ _13999_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23840_ _10090_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__clkbuf_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35826_ clknet_leaf_380_CLK _03940_ VGND VGND VPWR VPWR registers\[8\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35757_ clknet_leaf_389_CLK _03871_ VGND VGND VPWR VPWR registers\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_23771_ _10053_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32969_ clknet_leaf_193_CLK _01083_ VGND VGND VPWR VPWR registers\[53\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20983_ _07303_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__buf_6
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_509 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25510_ registers\[4\]\[21\] _10349_ _11034_ VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__mux2_1
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22722_ _09359_ _09362_ _09116_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__o21ba_1
X_34708_ clknet_leaf_94_CLK _02822_ VGND VGND VPWR VPWR registers\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_26490_ _11553_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35688_ clknet_leaf_459_CLK _03802_ VGND VGND VPWR VPWR registers\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25441_ _10997_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34639_ clknet_leaf_118_CLK _02753_ VGND VGND VPWR VPWR registers\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_22653_ registers\[4\]\[56\] registers\[5\]\[56\] registers\[6\]\[56\] registers\[7\]\[56\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__mux4_1
XFILLER_213_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21604_ _08271_ _08276_ _08073_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__o21ba_1
X_28160_ _12464_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__clkbuf_1
X_25372_ _10961_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22584_ registers\[52\]\[54\] registers\[53\]\[54\] registers\[54\]\[54\] registers\[55\]\[54\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__mux4_1
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27111_ _11818_ registers\[38\]\[42\] _11909_ VGND VGND VPWR VPWR _11912_ sky130_fd_sc_hd__mux2_1
X_24323_ net18 VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__clkbuf_4
X_28091_ _11851_ registers\[31\]\[58\] _12419_ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__mux2_1
X_21535_ _07347_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__buf_6
XFILLER_182_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27042_ _11875_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24254_ _10310_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21466_ registers\[4\]\[22\] registers\[5\]\[22\] registers\[6\]\[22\] registers\[7\]\[22\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__mux4_1
XFILLER_107_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23205_ _09733_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
X_20417_ registers\[16\]\[58\] registers\[17\]\[58\] registers\[18\]\[58\] registers\[19\]\[58\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__mux4_1
X_24185_ _10272_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
X_21397_ registers\[24\]\[20\] registers\[25\]\[20\] registers\[26\]\[20\] registers\[27\]\[20\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__mux4_1
XFILLER_218_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23136_ net8 VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__buf_6
X_20348_ _07051_ _07054_ _06855_ _06856_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__o211a_1
XFILLER_190_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28993_ _12902_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__clkbuf_1
XTAP_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27944_ registers\[32\]\[52\] _10414_ _12348_ VGND VGND VPWR VPWR _12351_ sky130_fd_sc_hd__mux2_1
XTAP_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23067_ _09641_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
XTAP_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20279_ registers\[56\]\[54\] registers\[57\]\[54\] registers\[58\]\[54\] registers\[59\]\[54\]
+ _06987_ _06777_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__mux4_1
XTAP_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22018_ registers\[60\]\[38\] registers\[61\]\[38\] registers\[62\]\[38\] registers\[63\]\[38\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__mux4_1
XFILLER_88_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27875_ _12314_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__clkbuf_1
XTAP_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29614_ _13260_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__clkbuf_1
X_26826_ net12 VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__clkbuf_4
XTAP_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29545_ _13224_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__clkbuf_1
X_23969_ _10157_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
X_26757_ registers\[40\]\[33\] _10374_ _11691_ VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__mux2_1
XFILLER_91_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16510_ registers\[0\]\[12\] registers\[1\]\[12\] registers\[2\]\[12\] registers\[3\]\[12\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15012_ sky130_fd_sc_hd__mux4_1
X_25708_ _11085_ VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__clkbuf_8
X_26688_ registers\[40\]\[0\] _10303_ _11658_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__mux2_1
X_17490_ _14555_ VGND VGND VPWR VPWR _15964_ sky130_fd_sc_hd__clkbuf_4
X_29476_ _09782_ registers\[21\]\[43\] _13184_ VGND VGND VPWR VPWR _13188_ sky130_fd_sc_hd__mux2_1
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16441_ _14584_ VGND VGND VPWR VPWR _14945_ sky130_fd_sc_hd__buf_2
X_28427_ _11782_ registers\[28\]\[25\] _12599_ VGND VGND VPWR VPWR _12605_ sky130_fd_sc_hd__mux2_1
X_25639_ registers\[48\]\[17\] _10340_ _11097_ VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__mux2_1
XFILLER_231_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ _14872_ _14877_ _14585_ VGND VGND VPWR VPWR _14878_ sky130_fd_sc_hd__o21ba_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19160_ _05755_ _05899_ _05900_ _05759_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__a22o_1
X_28358_ _12568_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18111_ _14491_ _04878_ _04879_ _14501_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a22o_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27309_ registers\[36\]\[8\] _10321_ _12007_ VGND VGND VPWR VPWR _12016_ sky130_fd_sc_hd__mux2_1
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ registers\[12\]\[20\] registers\[13\]\[20\] registers\[14\]\[20\] registers\[15\]\[20\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__mux4_1
X_28289_ _12532_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30320_ _13631_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__clkbuf_1
X_18042_ registers\[56\]\[56\] registers\[57\]\[56\] registers\[58\]\[56\] registers\[59\]\[56\]
+ _04751_ _04541_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__mux4_1
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30251_ _13595_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30182_ registers\[16\]\[58\] _13056_ _13550_ VGND VGND VPWR VPWR _13559_ sky130_fd_sc_hd__mux2_1
X_19993_ _06433_ _06708_ _06709_ _06439_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__a22o_1
XFILLER_99_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18944_ _05116_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__clkbuf_4
X_34990_ clknet_leaf_394_CLK _03104_ VGND VGND VPWR VPWR registers\[21\]\[32\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1420 _00182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1431 _05008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1442 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33941_ clknet_leaf_117_CLK _02055_ VGND VGND VPWR VPWR registers\[37\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18875_ registers\[8\]\[14\] registers\[9\]\[14\] registers\[10\]\[14\] registers\[11\]\[14\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__mux4_1
XFILLER_80_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1453 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1464 _05159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1475 _05476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1486 _07289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17826_ registers\[40\]\[50\] registers\[41\]\[50\] registers\[42\]\[50\] registers\[43\]\[50\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__mux4_1
XANTENNA_1497 _07326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33872_ clknet_leaf_127_CLK _01986_ VGND VGND VPWR VPWR registers\[38\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35611_ clknet_leaf_16_CLK _03725_ VGND VGND VPWR VPWR registers\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_32823_ clknet_leaf_330_CLK _00937_ VGND VGND VPWR VPWR registers\[55\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_17757_ registers\[44\]\[48\] registers\[45\]\[48\] registers\[46\]\[48\] registers\[47\]\[48\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__mux4_1
XFILLER_242_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35542_ clknet_leaf_82_CLK _03656_ VGND VGND VPWR VPWR registers\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_16708_ _14500_ VGND VGND VPWR VPWR _15204_ sky130_fd_sc_hd__clkbuf_4
X_32754_ clknet_leaf_363_CLK _00868_ VGND VGND VPWR VPWR registers\[56\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17688_ registers\[36\]\[46\] registers\[37\]\[46\] registers\[38\]\[46\] registers\[39\]\[46\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__mux4_1
X_31705_ registers\[59\]\[11\] net3 _14359_ VGND VGND VPWR VPWR _14361_ sky130_fd_sc_hd__mux2_1
XFILLER_39_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19427_ _05890_ _06158_ _06159_ _05893_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__a22o_1
X_35473_ clknet_leaf_76_CLK _03587_ VGND VGND VPWR VPWR registers\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16639_ _14863_ _15133_ _15136_ _14867_ VGND VGND VPWR VPWR _15137_ sky130_fd_sc_hd__a22o_1
X_32685_ clknet_leaf_372_CLK _00799_ VGND VGND VPWR VPWR registers\[57\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34424_ clknet_leaf_309_CLK _02538_ VGND VGND VPWR VPWR registers\[30\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_31636_ _14324_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__clkbuf_1
X_19358_ _05090_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__buf_6
XFILLER_91_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_241_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18309_ _05060_ _05063_ _05066_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a22o_1
XFILLER_176_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34355_ clknet_leaf_413_CLK _02469_ VGND VGND VPWR VPWR registers\[31\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31567_ _14276_ VGND VGND VPWR VPWR _14288_ sky130_fd_sc_hd__buf_6
X_19289_ _05095_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__buf_8
XFILLER_164_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33306_ clknet_leaf_31_CLK _01420_ VGND VGND VPWR VPWR registers\[47\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_21320_ registers\[12\]\[18\] registers\[13\]\[18\] registers\[14\]\[18\] registers\[15\]\[18\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__mux4_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30518_ _13736_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34286_ clknet_leaf_352_CLK _02400_ VGND VGND VPWR VPWR registers\[32\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31498_ _09778_ registers\[6\]\[41\] _14250_ VGND VGND VPWR VPWR _14252_ sky130_fd_sc_hd__mux2_1
X_36025_ clknet_leaf_332_CLK _04139_ VGND VGND VPWR VPWR registers\[63\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_33237_ clknet_leaf_70_CLK _01351_ VGND VGND VPWR VPWR registers\[48\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_21251_ _07928_ _07933_ _07730_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__o21ba_2
X_30449_ _09810_ registers\[14\]\[56\] _13693_ VGND VGND VPWR VPWR _13700_ sky130_fd_sc_hd__mux2_1
XFILLER_239_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20202_ _05042_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__buf_8
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33168_ clknet_leaf_139_CLK _01282_ VGND VGND VPWR VPWR registers\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21182_ _07347_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__buf_6
XFILLER_137_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20133_ _06576_ _06844_ _06845_ _06579_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__a22o_1
X_32119_ clknet_leaf_465_CLK _00035_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dfxtp_1
X_25990_ _11290_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
X_33099_ clknet_leaf_164_CLK _01213_ VGND VGND VPWR VPWR registers\[51\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20064_ _05090_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__buf_4
XFILLER_135_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24941_ _10703_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24872_ _09531_ registers\[53\]\[8\] _10658_ VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__mux2_1
X_27660_ _12201_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23823_ _10080_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__clkbuf_1
X_26611_ _11617_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__clkbuf_1
X_35809_ clknet_leaf_483_CLK _03923_ VGND VGND VPWR VPWR registers\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_27591_ _12165_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__clkbuf_1
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26542_ _11580_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_317 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29330_ _09771_ registers\[22\]\[38\] _13102_ VGND VGND VPWR VPWR _13111_ sky130_fd_sc_hd__mux2_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23754_ _10044_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_339 _00089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20966_ _07581_ _07655_ _07656_ _07584_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__a22o_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22705_ registers\[60\]\[58\] registers\[61\]\[58\] registers\[62\]\[58\] registers\[63\]\[58\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__mux4_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29261_ _09668_ registers\[22\]\[5\] _13069_ VGND VGND VPWR VPWR _13075_ sky130_fd_sc_hd__mux2_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26473_ _11544_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__clkbuf_1
X_23685_ _10006_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20897_ _07586_ _07587_ _07588_ _07589_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__a22o_1
XFILLER_198_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28212_ _11837_ registers\[30\]\[51\] _12490_ VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__mux2_1
X_25424_ _10988_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22636_ registers\[32\]\[56\] registers\[33\]\[56\] registers\[34\]\[56\] registers\[35\]\[56\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__mux4_1
X_29192_ registers\[23\]\[45\] _13029_ _13019_ VGND VGND VPWR VPWR _13030_ sky130_fd_sc_hd__mux2_1
XFILLER_167_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25355_ _10952_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_1
X_28143_ _12455_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__clkbuf_1
X_22567_ _09109_ _09211_ _09212_ _09114_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__a22o_1
XFILLER_167_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24306_ _10345_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
X_28074_ _12363_ VGND VGND VPWR VPWR _12419_ sky130_fd_sc_hd__buf_4
X_21518_ _08189_ _08192_ _08054_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__o21ba_1
XFILLER_194_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25286_ _10915_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_1
X_22498_ _09142_ _09145_ _09116_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__o21ba_1
XFILLER_186_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27025_ _11732_ registers\[38\]\[1\] _11865_ VGND VGND VPWR VPWR _11867_ sky130_fd_sc_hd__mux2_1
XFILLER_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24237_ _10299_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21449_ _07324_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__buf_4
XFILLER_5_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24168_ _10263_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_857 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23119_ registers\[39\]\[10\] _09678_ _09679_ VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__mux2_1
X_24099_ _10226_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
X_28976_ _12893_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__clkbuf_1
X_16990_ _14548_ VGND VGND VPWR VPWR _15478_ sky130_fd_sc_hd__buf_6
XFILLER_7_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27927_ registers\[32\]\[44\] _10397_ _12337_ VGND VGND VPWR VPWR _12342_ sky130_fd_sc_hd__mux2_1
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ registers\[52\]\[8\] registers\[53\]\[8\] registers\[54\]\[8\] registers\[55\]\[8\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__mux4_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27858_ registers\[32\]\[11\] _10328_ _12304_ VGND VGND VPWR VPWR _12306_ sky130_fd_sc_hd__mux2_1
XFILLER_23_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17611_ _04289_ _04393_ _04394_ _04292_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a22o_1
XFILLER_114_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26809_ registers\[40\]\[58\] _10426_ _11713_ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__mux2_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18591_ _05116_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__buf_4
XFILLER_188_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27789_ _12269_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29528_ _13215_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__clkbuf_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ registers\[28\]\[41\] registers\[29\]\[41\] registers\[30\]\[41\] registers\[31\]\[41\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__mux4_1
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_840 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_851 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_862 _09306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29459_ _09764_ registers\[21\]\[35\] _13173_ VGND VGND VPWR VPWR _13179_ sky130_fd_sc_hd__mux2_1
X_17473_ registers\[40\]\[40\] registers\[41\]\[40\] registers\[42\]\[40\] registers\[43\]\[40\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15947_ sky130_fd_sc_hd__mux4_1
XFILLER_229_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_873 _09514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_229_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_884 _09580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_895 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19212_ registers\[40\]\[24\] registers\[41\]\[24\] registers\[42\]\[24\] registers\[43\]\[24\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__mux4_1
X_16424_ registers\[56\]\[10\] registers\[57\]\[10\] registers\[58\]\[10\] registers\[59\]\[10\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _14928_ sky130_fd_sc_hd__mux4_1
X_32470_ clknet_leaf_62_CLK _00584_ VGND VGND VPWR VPWR registers\[60\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31421_ _14211_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__clkbuf_1
X_19143_ _05042_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__buf_4
X_16355_ _14500_ VGND VGND VPWR VPWR _14861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_146_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34140_ clknet_leaf_22_CLK _02254_ VGND VGND VPWR VPWR registers\[34\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_16286_ _14540_ _14790_ _14793_ _14551_ VGND VGND VPWR VPWR _14794_ sky130_fd_sc_hd__a22o_1
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31352_ registers\[7\]\[36\] net30 _14168_ VGND VGND VPWR VPWR _14175_ sky130_fd_sc_hd__mux2_1
X_19074_ _05547_ _05815_ _05816_ _05550_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a22o_1
XFILLER_172_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30303_ registers\[15\]\[51\] _13042_ _13621_ VGND VGND VPWR VPWR _13623_ sky130_fd_sc_hd__mux2_1
X_18025_ _04793_ _04796_ _04630_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__o21ba_1
XFILLER_199_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34071_ clknet_leaf_109_CLK _02185_ VGND VGND VPWR VPWR registers\[35\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_31283_ registers\[7\]\[3\] net34 _14135_ VGND VGND VPWR VPWR _14139_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33022_ clknet_leaf_268_CLK _01136_ VGND VGND VPWR VPWR registers\[52\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30234_ _13586_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30165_ _13494_ VGND VGND VPWR VPWR _13550_ sky130_fd_sc_hd__buf_4
X_19976_ registers\[16\]\[45\] registers\[17\]\[45\] registers\[18\]\[45\] registers\[19\]\[45\]
+ _06386_ _06387_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux4_1
XFILLER_45_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18927_ _05540_ _05672_ _05673_ _05545_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__a22o_1
XFILLER_132_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34973_ clknet_leaf_491_CLK _03087_ VGND VGND VPWR VPWR registers\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_30096_ registers\[16\]\[17\] _12970_ _13506_ VGND VGND VPWR VPWR _13514_ sky130_fd_sc_hd__mux2_1
XANTENNA_1250 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1261 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33924_ clknet_leaf_253_CLK _02038_ VGND VGND VPWR VPWR registers\[38\]\[54\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1272 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1283 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18858_ _05607_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1294 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17809_ _04583_ _04586_ _15963_ _15964_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__o211a_1
X_33855_ clknet_leaf_296_CLK _01969_ VGND VGND VPWR VPWR registers\[3\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18789_ _05076_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__clkbuf_4
X_20820_ _07325_ _07513_ _07514_ _07336_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__a22o_1
X_32806_ clknet_leaf_437_CLK _00920_ VGND VGND VPWR VPWR registers\[55\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33786_ clknet_leaf_280_CLK _01900_ VGND VGND VPWR VPWR registers\[40\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_30998_ _13988_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1062 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35525_ clknet_leaf_230_CLK _03639_ VGND VGND VPWR VPWR registers\[13\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20751_ _07313_ _07446_ _07447_ _07322_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a22o_1
X_32737_ clknet_leaf_44_CLK _00851_ VGND VGND VPWR VPWR registers\[56\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35456_ clknet_leaf_239_CLK _03570_ VGND VGND VPWR VPWR registers\[14\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23470_ _09556_ registers\[19\]\[20\] _09892_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__mux2_1
XFILLER_51_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20682_ registers\[16\]\[0\] registers\[17\]\[0\] registers\[18\]\[0\] registers\[19\]\[0\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__mux4_1
X_32668_ clknet_leaf_39_CLK _00782_ VGND VGND VPWR VPWR registers\[57\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22421_ registers\[20\]\[49\] registers\[21\]\[49\] registers\[22\]\[49\] registers\[23\]\[49\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__mux4_1
X_34407_ clknet_leaf_455_CLK _02521_ VGND VGND VPWR VPWR registers\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_31619_ _14315_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35387_ clknet_leaf_304_CLK _03501_ VGND VGND VPWR VPWR registers\[15\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_32599_ clknet_leaf_65_CLK _00713_ VGND VGND VPWR VPWR registers\[58\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25140_ net43 VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__buf_2
X_22352_ _08982_ _08989_ _08996_ _09003_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__or4_4
XFILLER_17_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34338_ clknet_leaf_470_CLK _02452_ VGND VGND VPWR VPWR registers\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21303_ _07316_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__clkbuf_4
XFILLER_191_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25071_ _10784_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
X_22283_ _08936_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_2
X_34269_ clknet_leaf_20_CLK _02383_ VGND VGND VPWR VPWR registers\[32\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24022_ _10186_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
X_36008_ clknet_leaf_436_CLK _04122_ VGND VGND VPWR VPWR registers\[63\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_21234_ _07640_ _07915_ _07916_ _07646_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__a22o_1
XFILLER_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28830_ _11780_ registers\[25\]\[24\] _12812_ VGND VGND VPWR VPWR _12817_ sky130_fd_sc_hd__mux2_1
X_21165_ _07846_ _07849_ _07711_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20116_ _06826_ _06829_ _06523_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o21ba_1
X_28761_ _12780_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__clkbuf_1
X_25973_ _11281_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
X_21096_ _07324_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27712_ registers\[33\]\[6\] _10317_ _12222_ VGND VGND VPWR VPWR _12229_ sky130_fd_sc_hd__mux2_1
XFILLER_63_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20047_ _06525_ _06761_ _06762_ _06528_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__a22o_1
X_24924_ _10694_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28692_ _12744_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27643_ _12192_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__clkbuf_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24855_ _10657_ VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__buf_4
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_103 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23806_ _10071_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27574_ _12156_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__clkbuf_1
X_24786_ _09580_ registers\[54\]\[31\] _10620_ VGND VGND VPWR VPWR _10622_ sky130_fd_sc_hd__mux2_1
XANTENNA_125 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _08656_ _08659_ _08430_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__o21ba_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29313_ _13068_ VGND VGND VPWR VPWR _13102_ sky130_fd_sc_hd__buf_4
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26525_ _10840_ registers\[42\]\[52\] _11569_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__mux2_1
X_23737_ _10035_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_158 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_169 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20949_ _07312_ VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__clkbuf_4
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29244_ registers\[23\]\[62\] _13064_ _12934_ VGND VGND VPWR VPWR _13065_ sky130_fd_sc_hd__mux2_1
XFILLER_198_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23668_ _09997_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_1
X_26456_ _11535_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22619_ registers\[8\]\[55\] registers\[9\]\[55\] registers\[10\]\[55\] registers\[11\]\[55\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__mux4_2
X_25407_ _10979_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_1
X_26387_ _11499_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29175_ net35 VGND VGND VPWR VPWR _13018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23599_ _09961_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
X_16140_ registers\[32\]\[2\] registers\[33\]\[2\] registers\[34\]\[2\] registers\[35\]\[2\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14652_ sky130_fd_sc_hd__mux4_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25338_ _10943_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__clkbuf_1
X_28126_ _11750_ registers\[30\]\[10\] _12446_ VGND VGND VPWR VPWR _12447_ sky130_fd_sc_hd__mux2_1
XFILLER_155_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16071_ _14584_ VGND VGND VPWR VPWR _14585_ sky130_fd_sc_hd__buf_2
XFILLER_108_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25269_ _10906_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__clkbuf_1
X_28057_ _12410_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27008_ net57 VGND VGND VPWR VPWR _11855_ sky130_fd_sc_hd__buf_2
XFILLER_108_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19830_ _06441_ _06550_ _06551_ _06445_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a22o_1
XFILLER_155_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19761_ registers\[4\]\[39\] registers\[5\]\[39\] registers\[6\]\[39\] registers\[7\]\[39\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__mux4_1
X_16973_ registers\[20\]\[25\] registers\[21\]\[25\] registers\[22\]\[25\] registers\[23\]\[25\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15462_ sky130_fd_sc_hd__mux4_1
X_28959_ registers\[24\]\[21\] _10349_ _12883_ VGND VGND VPWR VPWR _12885_ sky130_fd_sc_hd__mux2_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18712_ _05444_ _05451_ _05458_ _05465_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__or4_4
XFILLER_209_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31970_ clknet_leaf_5_CLK _00140_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_1
X_19692_ registers\[24\]\[37\] registers\[25\]\[37\] registers\[26\]\[37\] registers\[27\]\[37\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__mux4_1
XFILLER_232_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 DW[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_6
X_18643_ registers\[32\]\[8\] registers\[33\]\[8\] registers\[34\]\[8\] registers\[35\]\[8\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__mux4_1
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30921_ _13948_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33640_ clknet_leaf_430_CLK _01754_ VGND VGND VPWR VPWR registers\[42\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_30852_ _09808_ registers\[11\]\[55\] _13906_ VGND VGND VPWR VPWR _13912_ sky130_fd_sc_hd__mux2_1
X_18574_ _05197_ _05329_ _05330_ _05202_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__a22o_1
XFILLER_149_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17525_ registers\[56\]\[41\] registers\[57\]\[41\] registers\[58\]\[41\] registers\[59\]\[41\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__mux4_1
X_33571_ clknet_leaf_57_CLK _01685_ VGND VGND VPWR VPWR registers\[43\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_30783_ _09717_ registers\[11\]\[22\] _13873_ VGND VGND VPWR VPWR _13876_ sky130_fd_sc_hd__mux2_1
XANTENNA_670 _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35310_ clknet_leaf_397_CLK _03424_ VGND VGND VPWR VPWR registers\[16\]\[32\] sky130_fd_sc_hd__dfxtp_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32522_ clknet_leaf_178_CLK _00636_ VGND VGND VPWR VPWR registers\[60\]\[60\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_681 _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_692 _06823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17456_ _15927_ _15930_ _15620_ _15621_ VGND VGND VPWR VPWR _15931_ sky130_fd_sc_hd__o211a_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_978 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16407_ _14588_ _14910_ _14911_ _14598_ VGND VGND VPWR VPWR _14912_ sky130_fd_sc_hd__a22o_1
X_35241_ clknet_leaf_404_CLK _03355_ VGND VGND VPWR VPWR registers\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32453_ clknet_leaf_213_CLK _00567_ VGND VGND VPWR VPWR registers\[29\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17387_ _15825_ _15862_ _15863_ _15828_ VGND VGND VPWR VPWR _15864_ sky130_fd_sc_hd__a22o_1
XFILLER_220_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31404_ registers\[7\]\[61\] net58 _14134_ VGND VGND VPWR VPWR _14202_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19126_ registers\[8\]\[21\] registers\[9\]\[21\] registers\[10\]\[21\] registers\[11\]\[21\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__mux4_1
XFILLER_158_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16338_ _14601_ _14843_ _14844_ _14611_ VGND VGND VPWR VPWR _14845_ sky130_fd_sc_hd__a22o_1
XFILLER_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35172_ clknet_leaf_447_CLK _03286_ VGND VGND VPWR VPWR registers\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_32384_ clknet_leaf_293_CLK _00498_ VGND VGND VPWR VPWR registers\[61\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34123_ clknet_leaf_157_CLK _02237_ VGND VGND VPWR VPWR registers\[35\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31335_ registers\[7\]\[28\] net21 _14157_ VGND VGND VPWR VPWR _14166_ sky130_fd_sc_hd__mux2_1
X_19057_ _05797_ _05800_ _05494_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__o21ba_1
X_16269_ _14774_ _14777_ _14614_ VGND VGND VPWR VPWR _14778_ sky130_fd_sc_hd__o21ba_1
X_18008_ registers\[44\]\[55\] registers\[45\]\[55\] registers\[46\]\[55\] registers\[47\]\[55\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__mux4_1
XFILLER_195_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34054_ clknet_leaf_261_CLK _02168_ VGND VGND VPWR VPWR registers\[36\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_31266_ _14129_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33005_ clknet_leaf_373_CLK _01119_ VGND VGND VPWR VPWR registers\[52\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_30217_ registers\[15\]\[10\] _12955_ _13577_ VGND VGND VPWR VPWR _13578_ sky130_fd_sc_hd__mux2_1
XFILLER_113_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31197_ _14093_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ registers\[56\]\[45\] registers\[57\]\[45\] registers\[58\]\[45\] registers\[59\]\[45\]
+ _06644_ _06434_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__mux4_1
X_30148_ _13541_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34956_ clknet_leaf_141_CLK _03070_ VGND VGND VPWR VPWR registers\[22\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22970_ _09575_ registers\[62\]\[29\] _09557_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__mux2_1
XANTENNA_1080 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_228_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30079_ registers\[16\]\[9\] _12953_ _13495_ VGND VGND VPWR VPWR _13505_ sky130_fd_sc_hd__mux2_1
XFILLER_56_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1091 _14520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21921_ _08581_ _08584_ _08416_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__o21ba_1
X_33907_ clknet_leaf_349_CLK _02021_ VGND VGND VPWR VPWR registers\[38\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_34887_ clknet_leaf_206_CLK _03001_ VGND VGND VPWR VPWR registers\[23\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_24640_ _09571_ registers\[55\]\[27\] _10536_ VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__mux2_1
XFILLER_167_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33838_ clknet_leaf_389_CLK _01952_ VGND VGND VPWR VPWR registers\[3\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_21852_ registers\[12\]\[33\] registers\[13\]\[33\] registers\[14\]\[33\] registers\[15\]\[33\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__mux4_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20803_ _07495_ _07498_ _07399_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__o21ba_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24571_ _09640_ registers\[56\]\[60\] _10439_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__mux2_1
X_21783_ registers\[4\]\[31\] registers\[5\]\[31\] registers\[6\]\[31\] registers\[7\]\[31\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__mux4_1
X_33769_ clknet_leaf_427_CLK _01883_ VGND VGND VPWR VPWR registers\[40\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23522_ _09609_ registers\[19\]\[45\] _09914_ VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__mux2_1
X_26310_ _10760_ registers\[43\]\[14\] _11454_ VGND VGND VPWR VPWR _11459_ sky130_fd_sc_hd__mux2_1
X_20734_ _07410_ _07417_ _07424_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__or4_4
X_27290_ _12005_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__clkbuf_1
X_35508_ clknet_leaf_416_CLK _03622_ VGND VGND VPWR VPWR registers\[13\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26241_ _11422_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35439_ clknet_leaf_375_CLK _03553_ VGND VGND VPWR VPWR registers\[14\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_23453_ _09540_ registers\[19\]\[12\] _09881_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__mux2_1
X_20665_ _07363_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22404_ registers\[48\]\[49\] registers\[49\]\[49\] registers\[50\]\[49\] registers\[51\]\[49\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__mux4_1
X_26172_ _11386_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23384_ registers\[39\]\[45\] _09786_ _09840_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__mux2_1
X_20596_ _07294_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__buf_12
XFILLER_176_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25123_ _10819_ registers\[52\]\[42\] _10815_ VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__mux2_1
X_22335_ registers\[52\]\[47\] registers\[53\]\[47\] registers\[54\]\[47\] registers\[55\]\[47\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__mux4_1
XFILLER_178_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29931_ _13427_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__clkbuf_1
X_25054_ _10730_ VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__buf_4
X_22266_ _07287_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__buf_6
XFILLER_136_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24005_ _10177_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
X_21217_ registers\[16\]\[15\] registers\[17\]\[15\] registers\[18\]\[15\] registers\[19\]\[15\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__mux4_1
XFILLER_105_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29862_ registers\[18\]\[34\] _13006_ _13386_ VGND VGND VPWR VPWR _13391_ sky130_fd_sc_hd__mux2_1
X_22197_ registers\[52\]\[43\] registers\[53\]\[43\] registers\[54\]\[43\] registers\[55\]\[43\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__mux4_1
XFILLER_105_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28813_ _11763_ registers\[25\]\[16\] _12801_ VGND VGND VPWR VPWR _12808_ sky130_fd_sc_hd__mux2_1
XFILLER_152_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21148_ _07586_ _07832_ _07833_ _07589_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__a22o_1
X_29793_ registers\[18\]\[1\] _12937_ _13353_ VGND VGND VPWR VPWR _13355_ sky130_fd_sc_hd__mux2_1
XFILLER_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28744_ _12771_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__clkbuf_1
X_21079_ _07763_ _07766_ _07730_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__o21ba_2
X_25956_ _11272_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24907_ _10685_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28675_ _12735_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__clkbuf_1
X_25887_ _11236_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27626_ _12183_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__clkbuf_1
X_24838_ _09632_ registers\[54\]\[56\] _10642_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__mux2_1
XFILLER_132_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27557_ _11859_ registers\[35\]\[62\] _12077_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__mux2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _09563_ registers\[54\]\[23\] _10609_ VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__mux2_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17310_ registers\[52\]\[35\] registers\[53\]\[35\] registers\[54\]\[35\] registers\[55\]\[35\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15789_ sky130_fd_sc_hd__mux4_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26508_ _10823_ registers\[42\]\[44\] _11558_ VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__mux2_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _05044_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__buf_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27488_ _11790_ registers\[35\]\[29\] _12100_ VGND VGND VPWR VPWR _12110_ sky130_fd_sc_hd__mux2_1
XFILLER_202_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29227_ _13053_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17241_ registers\[48\]\[33\] registers\[49\]\[33\] registers\[50\]\[33\] registers\[51\]\[33\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15722_ sky130_fd_sc_hd__mux4_1
XFILLER_35_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26439_ _10754_ registers\[42\]\[11\] _11525_ VGND VGND VPWR VPWR _11527_ sky130_fd_sc_hd__mux2_1
XFILLER_74_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17172_ registers\[56\]\[31\] registers\[57\]\[31\] registers\[58\]\[31\] registers\[59\]\[31\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15655_ sky130_fd_sc_hd__mux4_1
X_29158_ registers\[23\]\[34\] _13006_ _12998_ VGND VGND VPWR VPWR _13007_ sky130_fd_sc_hd__mux2_1
XFILLER_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16123_ registers\[12\]\[1\] registers\[13\]\[1\] registers\[14\]\[1\] registers\[15\]\[1\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _14636_ sky130_fd_sc_hd__mux4_1
X_28109_ _11734_ registers\[30\]\[2\] _12435_ VGND VGND VPWR VPWR _12438_ sky130_fd_sc_hd__mux2_1
XFILLER_122_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29089_ net4 VGND VGND VPWR VPWR _12960_ sky130_fd_sc_hd__buf_4
XFILLER_182_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31120_ registers\[0\]\[54\] _13048_ _14048_ VGND VGND VPWR VPWR _14053_ sky130_fd_sc_hd__mux2_1
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16054_ _14567_ VGND VGND VPWR VPWR _14568_ sky130_fd_sc_hd__buf_4
XFILLER_108_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31051_ registers\[0\]\[21\] _12979_ _14015_ VGND VGND VPWR VPWR _14017_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19813_ _06530_ _06531_ _06534_ _06535_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__a22o_1
X_30002_ _13464_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34810_ clknet_leaf_304_CLK _02924_ VGND VGND VPWR VPWR registers\[24\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19744_ registers\[32\]\[39\] registers\[33\]\[39\] registers\[34\]\[39\] registers\[35\]\[39\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__mux4_1
X_35790_ clknet_leaf_108_CLK _03904_ VGND VGND VPWR VPWR registers\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_16956_ registers\[60\]\[25\] registers\[61\]\[25\] registers\[62\]\[25\] registers\[63\]\[25\]
+ _15413_ _15207_ VGND VGND VPWR VPWR _15445_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34741_ clknet_leaf_413_CLK _02855_ VGND VGND VPWR VPWR registers\[25\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31953_ clknet_leaf_0_CLK _00161_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
X_19675_ registers\[36\]\[37\] registers\[37\]\[37\] registers\[38\]\[37\] registers\[39\]\[37\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__mux4_1
XFILLER_65_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16887_ registers\[56\]\[23\] registers\[57\]\[23\] registers\[58\]\[23\] registers\[59\]\[23\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15378_ sky130_fd_sc_hd__mux4_1
XFILLER_53_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18626_ registers\[8\]\[7\] registers\[9\]\[7\] registers\[10\]\[7\] registers\[11\]\[7\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__mux4_1
X_30904_ _13939_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__clkbuf_1
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34672_ clknet_leaf_411_CLK _02786_ VGND VGND VPWR VPWR registers\[26\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_31884_ _09758_ registers\[49\]\[32\] _14452_ VGND VGND VPWR VPWR _14455_ sky130_fd_sc_hd__mux2_1
XFILLER_92_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33623_ clknet_leaf_135_CLK _01737_ VGND VGND VPWR VPWR registers\[42\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_18557_ registers\[0\]\[5\] registers\[1\]\[5\] registers\[2\]\[5\] registers\[3\]\[5\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__mux4_1
X_30835_ _09791_ registers\[11\]\[47\] _13895_ VGND VGND VPWR VPWR _13903_ sky130_fd_sc_hd__mux2_1
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17508_ registers\[28\]\[40\] registers\[29\]\[40\] registers\[30\]\[40\] registers\[31\]\[40\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__mux4_1
X_33554_ clknet_leaf_125_CLK _01668_ VGND VGND VPWR VPWR registers\[43\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18488_ registers\[8\]\[3\] registers\[9\]\[3\] registers\[10\]\[3\] registers\[11\]\[3\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__mux4_1
X_30766_ _09687_ registers\[11\]\[14\] _13862_ VGND VGND VPWR VPWR _13867_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32505_ clknet_leaf_332_CLK _00619_ VGND VGND VPWR VPWR registers\[60\]\[43\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_14 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ _15883_ _15898_ _15907_ _15914_ VGND VGND VPWR VPWR _15915_ sky130_fd_sc_hd__or4_4
X_33485_ clknet_leaf_172_CLK _01599_ VGND VGND VPWR VPWR registers\[45\]\[63\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_25 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30697_ _13830_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_36 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_47 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35224_ clknet_leaf_7_CLK _03338_ VGND VGND VPWR VPWR registers\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_20450_ registers\[20\]\[59\] registers\[21\]\[59\] registers\[22\]\[59\] registers\[23\]\[59\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__mux4_1
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_58 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32436_ clknet_leaf_416_CLK _00550_ VGND VGND VPWR VPWR registers\[29\]\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_69 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_830 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19109_ _05843_ _05850_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__o21ba_1
X_35155_ clknet_leaf_102_CLK _03269_ VGND VGND VPWR VPWR registers\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20381_ _05040_ _07085_ _07086_ _05050_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__a22o_1
X_32367_ clknet_leaf_370_CLK _00481_ VGND VGND VPWR VPWR registers\[61\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34106_ clknet_leaf_281_CLK _02220_ VGND VGND VPWR VPWR registers\[35\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_22120_ _08462_ _08776_ _08777_ _08467_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__a22o_1
X_31318_ _14134_ VGND VGND VPWR VPWR _14157_ sky130_fd_sc_hd__buf_4
X_35086_ clknet_leaf_109_CLK _03200_ VGND VGND VPWR VPWR registers\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xoutput110 net110 VGND VGND VPWR VPWR D1[28] sky130_fd_sc_hd__buf_2
X_32298_ clknet_leaf_408_CLK _00412_ VGND VGND VPWR VPWR registers\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xoutput121 net121 VGND VGND VPWR VPWR D1[38] sky130_fd_sc_hd__buf_2
XFILLER_161_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput132 net132 VGND VGND VPWR VPWR D1[48] sky130_fd_sc_hd__buf_2
XFILLER_133_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput143 net143 VGND VGND VPWR VPWR D1[58] sky130_fd_sc_hd__buf_2
X_22051_ registers\[48\]\[39\] registers\[49\]\[39\] registers\[50\]\[39\] registers\[51\]\[39\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__mux4_1
X_34037_ clknet_leaf_343_CLK _02151_ VGND VGND VPWR VPWR registers\[36\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31249_ registers\[8\]\[51\] net47 _14119_ VGND VGND VPWR VPWR _14121_ sky130_fd_sc_hd__mux2_1
XTAP_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput154 net154 VGND VGND VPWR VPWR D2[0] sky130_fd_sc_hd__buf_2
Xoutput165 net165 VGND VGND VPWR VPWR D2[1] sky130_fd_sc_hd__buf_2
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21002_ registers\[4\]\[9\] registers\[5\]\[9\] registers\[6\]\[9\] registers\[7\]\[9\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__mux4_1
XFILLER_130_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput176 net176 VGND VGND VPWR VPWR D2[2] sky130_fd_sc_hd__buf_2
XFILLER_87_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput187 net187 VGND VGND VPWR VPWR D2[3] sky130_fd_sc_hd__buf_2
XTAP_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput198 net198 VGND VGND VPWR VPWR D2[4] sky130_fd_sc_hd__buf_2
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25810_ _10800_ registers\[47\]\[33\] _11192_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__mux2_1
XFILLER_29_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26790_ registers\[40\]\[49\] _10407_ _11702_ VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__mux2_1
X_35988_ clknet_leaf_63_CLK _04102_ VGND VGND VPWR VPWR registers\[63\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25741_ _10728_ registers\[47\]\[0\] _11159_ VGND VGND VPWR VPWR _11160_ sky130_fd_sc_hd__mux2_1
X_22953_ _09564_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
X_34939_ clknet_leaf_307_CLK _03053_ VGND VGND VPWR VPWR registers\[22\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_233_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21904_ _08469_ _08566_ _08567_ _08472_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a22o_1
X_28460_ _12622_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__clkbuf_1
X_22884_ _09517_ registers\[62\]\[1\] _09515_ VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__mux2_1
X_25672_ _11122_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27411_ _12069_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__clkbuf_1
X_21835_ _08462_ _08499_ _08500_ _08467_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__a22o_1
X_24623_ _09554_ registers\[55\]\[19\] _10525_ VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__mux2_1
XFILLER_231_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28391_ _11746_ registers\[28\]\[8\] _12577_ VGND VGND VPWR VPWR _12586_ sky130_fd_sc_hd__mux2_1
XFILLER_110_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24554_ _10497_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27342_ _12033_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_1
X_21766_ registers\[32\]\[31\] registers\[33\]\[31\] registers\[34\]\[31\] registers\[35\]\[31\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__mux4_1
XFILLER_212_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20717_ registers\[52\]\[1\] registers\[53\]\[1\] registers\[54\]\[1\] registers\[55\]\[1\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__mux4_1
X_23505_ _09592_ registers\[19\]\[37\] _09903_ VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__mux2_1
X_27273_ _11845_ registers\[37\]\[55\] _11991_ VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__mux2_1
XFILLER_180_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24485_ _09554_ registers\[56\]\[19\] _10451_ VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__mux2_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21697_ registers\[56\]\[29\] registers\[57\]\[29\] registers\[58\]\[29\] registers\[59\]\[29\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__mux4_1
X_29012_ _12912_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23436_ _09523_ registers\[19\]\[4\] _09870_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__mux2_1
X_26224_ _11413_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
X_20648_ _07314_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__buf_12
XFILLER_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26155_ _11377_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_192_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_192_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23367_ registers\[39\]\[37\] _09769_ _09829_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__mux2_1
X_20579_ _07277_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__buf_12
X_22318_ _08766_ _08969_ _08970_ _08771_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__a22o_1
XFILLER_139_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25106_ net31 VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__buf_2
XFILLER_164_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26086_ _10806_ registers\[45\]\[36\] _11334_ VGND VGND VPWR VPWR _11341_ sky130_fd_sc_hd__mux2_1
X_23298_ registers\[9\]\[48\] _09793_ _09776_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__mux2_1
XFILLER_30_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29914_ registers\[18\]\[59\] _13058_ _13408_ VGND VGND VPWR VPWR _13418_ sky130_fd_sc_hd__mux2_1
X_25037_ _10761_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
X_22249_ _08900_ _08903_ _08773_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29845_ registers\[18\]\[26\] _12989_ _13375_ VGND VGND VPWR VPWR _13382_ sky130_fd_sc_hd__mux2_1
XFILLER_239_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16810_ _15270_ _15279_ _15289_ _15303_ VGND VGND VPWR VPWR _15304_ sky130_fd_sc_hd__or4_4
X_29776_ _13345_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__clkbuf_1
X_17790_ _04294_ _04567_ _04568_ _04299_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a22o_1
XFILLER_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26988_ _11841_ registers\[3\]\[53\] _11835_ VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__mux2_1
XFILLER_232_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28727_ _12762_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__clkbuf_1
X_16741_ registers\[36\]\[19\] registers\[37\]\[19\] registers\[38\]\[19\] registers\[39\]\[19\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15236_ sky130_fd_sc_hd__mux4_1
XFILLER_143_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25939_ _10793_ registers\[46\]\[30\] _11263_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__mux2_1
XFILLER_235_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19460_ _06187_ _06188_ _06191_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__a22o_1
XFILLER_35_917 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28658_ _12726_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16672_ registers\[56\]\[17\] registers\[57\]\[17\] registers\[58\]\[17\] registers\[59\]\[17\]
+ _15066_ _14856_ VGND VGND VPWR VPWR _15169_ sky130_fd_sc_hd__mux4_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_6_25__f_CLK clknet_5_12_0_CLK VGND VGND VPWR VPWR clknet_6_25__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18411_ _05060_ _05169_ _05172_ _05066_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__a22o_1
XFILLER_185_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27609_ registers\[34\]\[21\] _10349_ _12173_ VGND VGND VPWR VPWR _12175_ sky130_fd_sc_hd__mux2_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ registers\[32\]\[29\] registers\[33\]\[29\] registers\[34\]\[29\] registers\[35\]\[29\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux4_1
XFILLER_222_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28589_ _11809_ registers\[27\]\[38\] _12681_ VGND VGND VPWR VPWR _12690_ sky130_fd_sc_hd__mux2_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30620_ registers\[12\]\[9\] _12953_ _13780_ VGND VGND VPWR VPWR _13790_ sky130_fd_sc_hd__mux2_1
X_18342_ _05104_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__buf_2
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _05015_ _05022_ _05029_ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__or4_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30551_ _09775_ registers\[13\]\[40\] _13753_ VGND VGND VPWR VPWR _13754_ sky130_fd_sc_hd__mux2_1
XFILLER_203_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17224_ _15633_ _15704_ _15705_ _15636_ VGND VGND VPWR VPWR _15706_ sky130_fd_sc_hd__a22o_1
X_33270_ clknet_leaf_336_CLK _01384_ VGND VGND VPWR VPWR registers\[48\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30482_ _13717_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 DW[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_8
XFILLER_11_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 DW[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_8
X_32221_ clknet_leaf_240_CLK _00335_ VGND VGND VPWR VPWR registers\[9\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput34 DW[3] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_8
XFILLER_128_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput45 DW[4] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_6
X_17155_ registers\[28\]\[30\] registers\[29\]\[30\] registers\[30\]\[30\] registers\[31\]\[30\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15639_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_183_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_183_CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput56 DW[5] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_6
Xinput67 R1[2] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_8
XFILLER_196_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput78 R3[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
X_16106_ _14491_ _14617_ _14618_ _14501_ VGND VGND VPWR VPWR _14619_ sky130_fd_sc_hd__a22o_1
Xinput89 WE VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_6
XFILLER_239_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32152_ clknet_leaf_31_CLK _00266_ VGND VGND VPWR VPWR registers\[39\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1006 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17086_ _15540_ _15555_ _15564_ _15571_ VGND VGND VPWR VPWR _15572_ sky130_fd_sc_hd__or4_4
XFILLER_143_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31103_ registers\[0\]\[46\] _13031_ _14037_ VGND VGND VPWR VPWR _14044_ sky130_fd_sc_hd__mux2_1
X_16037_ _14516_ VGND VGND VPWR VPWR _14551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32083_ clknet_leaf_490_CLK _00055_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35911_ clknet_leaf_210_CLK _04025_ VGND VGND VPWR VPWR registers\[7\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_31034_ registers\[0\]\[13\] _12962_ _14004_ VGND VGND VPWR VPWR _14008_ sky130_fd_sc_hd__mux2_1
XFILLER_135_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35842_ clknet_leaf_242_CLK _03956_ VGND VGND VPWR VPWR registers\[8\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_17988_ registers\[0\]\[54\] registers\[1\]\[54\] registers\[2\]\[54\] registers\[3\]\[54\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux4_1
X_19727_ _05125_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__buf_6
XFILLER_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16939_ _15290_ _15427_ _15428_ _15293_ VGND VGND VPWR VPWR _15429_ sky130_fd_sc_hd__a22o_1
X_35773_ clknet_leaf_288_CLK _03887_ VGND VGND VPWR VPWR registers\[0\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_32985_ clknet_leaf_67_CLK _01099_ VGND VGND VPWR VPWR registers\[52\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31936_ _09813_ registers\[49\]\[57\] _14474_ VGND VGND VPWR VPWR _14482_ sky130_fd_sc_hd__mux2_1
X_34724_ clknet_leaf_474_CLK _02838_ VGND VGND VPWR VPWR registers\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_19658_ registers\[24\]\[36\] registers\[25\]\[36\] registers\[26\]\[36\] registers\[27\]\[36\]
+ _06317_ _06318_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18609_ _05365_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
X_34655_ clknet_leaf_9_CLK _02769_ VGND VGND VPWR VPWR registers\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31867_ _09740_ registers\[49\]\[24\] _14441_ VGND VGND VPWR VPWR _14446_ sky130_fd_sc_hd__mux2_1
X_19589_ _05113_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__buf_4
XFILLER_225_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33606_ clknet_leaf_248_CLK _01720_ VGND VGND VPWR VPWR registers\[43\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_21620_ _07356_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__buf_6
X_30818_ _09773_ registers\[11\]\[39\] _13884_ VGND VGND VPWR VPWR _13894_ sky130_fd_sc_hd__mux2_1
X_34586_ clknet_leaf_20_CLK _02700_ VGND VGND VPWR VPWR registers\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_31798_ _14409_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33537_ clknet_leaf_257_CLK _01651_ VGND VGND VPWR VPWR registers\[44\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_21551_ _08126_ _08223_ _08224_ _08129_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__a22o_1
XFILLER_181_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30749_ _09670_ registers\[11\]\[6\] _13851_ VGND VGND VPWR VPWR _13858_ sky130_fd_sc_hd__mux2_1
XFILLER_194_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20502_ registers\[12\]\[61\] registers\[13\]\[61\] registers\[14\]\[61\] registers\[15\]\[61\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__mux4_1
XFILLER_21_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24270_ net63 VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__buf_4
XFILLER_166_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33468_ clknet_leaf_278_CLK _01582_ VGND VGND VPWR VPWR registers\[45\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_21482_ _08119_ _08156_ _08157_ _08124_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__a22o_1
XFILLER_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35207_ clknet_leaf_153_CLK _03321_ VGND VGND VPWR VPWR registers\[18\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23221_ registers\[9\]\[25\] _09742_ _09735_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__mux2_1
XFILLER_222_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20433_ registers\[48\]\[59\] registers\[49\]\[59\] registers\[50\]\[59\] registers\[51\]\[59\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__mux4_1
X_32419_ clknet_leaf_473_CLK _00533_ VGND VGND VPWR VPWR registers\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_174_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_174_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_36187_ clknet_leaf_93_CLK _00068_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
X_33399_ clknet_leaf_340_CLK _01513_ VGND VGND VPWR VPWR registers\[46\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35138_ clknet_leaf_241_CLK _03252_ VGND VGND VPWR VPWR registers\[1\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23152_ net14 VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__clkbuf_4
X_20364_ _07070_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__buf_4
XTAP_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22103_ registers\[24\]\[40\] registers\[25\]\[40\] registers\[26\]\[40\] registers\[27\]\[40\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__mux4_1
XTAP_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23083_ net83 net89 VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__nand2_8
X_27960_ registers\[32\]\[60\] _10430_ _12292_ VGND VGND VPWR VPWR _12359_ sky130_fd_sc_hd__mux2_1
XFILLER_162_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35069_ clknet_leaf_188_CLK _03183_ VGND VGND VPWR VPWR registers\[20\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_20295_ _05113_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__buf_4
XTAP_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26911_ _11789_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_1
X_22034_ _08418_ _08693_ _08694_ _08421_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__a22o_1
XTAP_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27891_ registers\[32\]\[27\] _10361_ _12315_ VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__mux2_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29630_ registers\[20\]\[52\] _13044_ _13266_ VGND VGND VPWR VPWR _13269_ sky130_fd_sc_hd__mux2_1
XTAP_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26842_ _11742_ registers\[3\]\[6\] _11730_ VGND VGND VPWR VPWR _11743_ sky130_fd_sc_hd__mux2_1
XTAP_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29561_ _13232_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26773_ _11703_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23985_ _09525_ registers\[5\]\[5\] _10161_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__mux2_1
XFILLER_68_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28512_ _11732_ registers\[27\]\[1\] _12648_ VGND VGND VPWR VPWR _12650_ sky130_fd_sc_hd__mux2_1
XFILLER_186_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25724_ _11149_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
X_29492_ _13196_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22936_ _09552_ registers\[62\]\[18\] _09536_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__mux2_1
X_28443_ _12613_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25655_ _11113_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22867_ registers\[16\]\[63\] registers\[17\]\[63\] registers\[18\]\[63\] registers\[19\]\[63\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__mux4_1
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24606_ _10526_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28374_ _12576_ VGND VGND VPWR VPWR _12577_ sky130_fd_sc_hd__buf_6
X_21818_ registers\[12\]\[32\] registers\[13\]\[32\] registers\[14\]\[32\] registers\[15\]\[32\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__mux4_1
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25586_ _11075_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
X_22798_ _09432_ _09435_ _07338_ _07340_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__o211a_1
XFILLER_244_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27325_ _12024_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkbuf_1
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24537_ _10488_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
X_21749_ _07372_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__clkbuf_4
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_936 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27256_ _11828_ registers\[37\]\[47\] _11980_ VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1058 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24468_ _10452_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26207_ _11404_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_165_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_165_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23419_ registers\[39\]\[62\] _09823_ _09657_ VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24399_ _10408_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
X_27187_ _11759_ registers\[37\]\[14\] _11947_ VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__mux2_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26138_ _10858_ registers\[45\]\[61\] _11300_ VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18960_ _05703_ _05706_ _05508_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26069_ _10789_ registers\[45\]\[28\] _11323_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__mux2_1
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17911_ _14516_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__buf_4
XANTENNA_1602 _14564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18891_ _05614_ _05623_ _05630_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__or4_2
XANTENNA_1613 _15508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1624 _15808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1635 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1646 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17842_ _14553_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29828_ registers\[18\]\[18\] _12972_ _13364_ VGND VGND VPWR VPWR _13373_ sky130_fd_sc_hd__mux2_1
XTAP_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1657 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1668 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1679 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17773_ _14515_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__buf_4
X_29759_ _13336_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19512_ registers\[52\]\[32\] registers\[53\]\[32\] registers\[54\]\[32\] registers\[55\]\[32\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux4_1
X_16724_ _15144_ _15216_ _15219_ _15147_ VGND VGND VPWR VPWR _15220_ sky130_fd_sc_hd__a22o_1
X_32770_ clknet_leaf_263_CLK _00884_ VGND VGND VPWR VPWR registers\[56\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_234_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19443_ _06031_ _06172_ _06175_ _06034_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__a22o_1
X_31721_ registers\[59\]\[19\] net11 _14359_ VGND VGND VPWR VPWR _14369_ sky130_fd_sc_hd__mux2_1
XFILLER_222_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16655_ registers\[16\]\[16\] registers\[17\]\[16\] registers\[18\]\[16\] registers\[19\]\[16\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15153_ sky130_fd_sc_hd__mux4_1
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34440_ clknet_leaf_212_CLK _02554_ VGND VGND VPWR VPWR registers\[30\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31652_ registers\[63\]\[50\] net46 _14332_ VGND VGND VPWR VPWR _14333_ sky130_fd_sc_hd__mux2_1
XFILLER_16_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19374_ _05125_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__buf_6
X_16586_ _14947_ _15084_ _15085_ _14950_ VGND VGND VPWR VPWR _15086_ sky130_fd_sc_hd__a22o_1
XFILLER_31_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30603_ _13781_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18325_ _05058_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__buf_12
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34371_ clknet_leaf_205_CLK _02485_ VGND VGND VPWR VPWR registers\[31\]\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31583_ _14296_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36110_ clknet_leaf_74_CLK _04224_ VGND VGND VPWR VPWR registers\[49\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_33322_ clknet_leaf_429_CLK _01436_ VGND VGND VPWR VPWR registers\[47\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_18256_ registers\[52\]\[63\] registers\[53\]\[63\] registers\[54\]\[63\] registers\[55\]\[63\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__mux4_1
X_30534_ _09758_ registers\[13\]\[32\] _13742_ VGND VGND VPWR VPWR _13745_ sky130_fd_sc_hd__mux2_1
XFILLER_31_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36041_ clknet_leaf_162_CLK _04155_ VGND VGND VPWR VPWR registers\[63\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17207_ _15683_ _15688_ _15612_ VGND VGND VPWR VPWR _15689_ sky130_fd_sc_hd__o21ba_1
X_33253_ clknet_leaf_439_CLK _01367_ VGND VGND VPWR VPWR registers\[48\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_30465_ _13636_ _10015_ VGND VGND VPWR VPWR _13708_ sky130_fd_sc_hd__nand2_8
Xclkbuf_leaf_156_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_156_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18187_ _04676_ _04951_ _04952_ _04681_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__a22o_1
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32204_ clknet_leaf_434_CLK _00318_ VGND VGND VPWR VPWR registers\[39\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17138_ _15616_ _15619_ _15620_ _15621_ VGND VGND VPWR VPWR _15622_ sky130_fd_sc_hd__o211a_1
XFILLER_190_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33184_ clknet_leaf_481_CLK _01298_ VGND VGND VPWR VPWR registers\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_30396_ _13672_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__clkbuf_1
X_32135_ clknet_leaf_460_CLK _00052_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17069_ _15548_ _15554_ _15277_ _15278_ VGND VGND VPWR VPWR _15555_ sky130_fd_sc_hd__o211a_1
XFILLER_98_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32066_ clknet_leaf_201_CLK _00244_ VGND VGND VPWR VPWR registers\[62\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_20080_ _05125_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__buf_6
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31017_ registers\[0\]\[5\] _12945_ _13993_ VGND VGND VPWR VPWR _13999_ sky130_fd_sc_hd__mux2_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35825_ clknet_leaf_381_CLK _03939_ VGND VGND VPWR VPWR registers\[8\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23770_ _09582_ registers\[29\]\[32\] _10050_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__mux2_1
X_20982_ registers\[40\]\[9\] registers\[41\]\[9\] registers\[42\]\[9\] registers\[43\]\[9\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__mux4_1
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32968_ clknet_leaf_191_CLK _01082_ VGND VGND VPWR VPWR registers\[53\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35756_ clknet_leaf_388_CLK _03870_ VGND VGND VPWR VPWR registers\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22721_ _09109_ _09360_ _09361_ _09114_ VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__a22o_1
X_34707_ clknet_leaf_104_CLK _02821_ VGND VGND VPWR VPWR registers\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_31919_ _09795_ registers\[49\]\[49\] _14463_ VGND VGND VPWR VPWR _14473_ sky130_fd_sc_hd__mux2_1
X_32899_ clknet_leaf_293_CLK _01013_ VGND VGND VPWR VPWR registers\[54\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35687_ clknet_leaf_460_CLK _03801_ VGND VGND VPWR VPWR registers\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22652_ registers\[12\]\[56\] registers\[13\]\[56\] registers\[14\]\[56\] registers\[15\]\[56\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__mux4_1
X_25440_ _10844_ registers\[50\]\[54\] _10992_ VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__mux2_1
X_34638_ clknet_leaf_118_CLK _02752_ VGND VGND VPWR VPWR registers\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21603_ _08272_ _08273_ _08274_ _08275_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__a22o_1
X_34569_ clknet_leaf_214_CLK _02683_ VGND VGND VPWR VPWR registers\[28\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_22583_ registers\[60\]\[54\] registers\[61\]\[54\] registers\[62\]\[54\] registers\[63\]\[54\]
+ _09227_ _09021_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_395_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_395_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25371_ _10775_ registers\[50\]\[21\] _10959_ VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__mux2_1
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27110_ _11911_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21534_ _08205_ _08208_ _08073_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__o21ba_1
X_24322_ _10356_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
X_28090_ _12427_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27041_ _11748_ registers\[38\]\[9\] _11865_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__mux2_1
XFILLER_182_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24253_ registers\[57\]\[2\] _10309_ _10305_ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_147_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_147_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21465_ registers\[12\]\[22\] registers\[13\]\[22\] registers\[14\]\[22\] registers\[15\]\[22\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__mux4_1
XFILLER_181_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23204_ registers\[9\]\[18\] _09695_ _09722_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__mux2_1
X_20416_ registers\[24\]\[58\] registers\[25\]\[58\] registers\[26\]\[58\] registers\[27\]\[58\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__mux4_1
XFILLER_107_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24184_ _09588_ registers\[58\]\[35\] _10266_ VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__mux2_1
X_21396_ _07372_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23135_ _09690_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
X_20347_ _06784_ _07052_ _07053_ _06788_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__a22o_1
XFILLER_49_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28992_ registers\[24\]\[37\] _10382_ _12894_ VGND VGND VPWR VPWR _12902_ sky130_fd_sc_hd__mux2_1
XFILLER_161_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27943_ _12350_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__clkbuf_1
X_23066_ _09640_ registers\[62\]\[60\] _09514_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__mux2_1
XFILLER_153_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20278_ _05078_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__buf_6
XTAP_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_752 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22017_ _07328_ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27874_ registers\[32\]\[19\] _10344_ _12304_ VGND VGND VPWR VPWR _12314_ sky130_fd_sc_hd__mux2_1
XFILLER_248_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29613_ registers\[20\]\[44\] _13027_ _13255_ VGND VGND VPWR VPWR _13260_ sky130_fd_sc_hd__mux2_1
XFILLER_114_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26825_ _11731_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__clkbuf_1
XTAP_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29544_ registers\[20\]\[11\] _12958_ _13222_ VGND VGND VPWR VPWR _13224_ sky130_fd_sc_hd__mux2_1
XFILLER_84_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26756_ _11694_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23968_ _09644_ registers\[60\]\[62\] _10088_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__mux2_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25707_ _11140_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29475_ _13187_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__clkbuf_1
X_22919_ _09541_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
X_26687_ _11657_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__buf_4
XFILLER_83_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23899_ _09575_ registers\[60\]\[29\] _10111_ VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__mux2_1
XFILLER_232_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28426_ _12604_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__clkbuf_1
X_16440_ _14801_ _14942_ _14943_ _14804_ VGND VGND VPWR VPWR _14944_ sky130_fd_sc_hd__a22o_1
X_25638_ _11104_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28357_ registers\[2\]\[56\] _10422_ _12561_ VGND VGND VPWR VPWR _12568_ sky130_fd_sc_hd__mux2_1
X_16371_ _14801_ _14873_ _14876_ _14804_ VGND VGND VPWR VPWR _14877_ sky130_fd_sc_hd__a22o_1
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25569_ _11066_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_386_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_386_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18110_ registers\[0\]\[58\] registers\[1\]\[58\] registers\[2\]\[58\] registers\[3\]\[58\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__mux4_1
X_27308_ _12015_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__clkbuf_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19090_ _05688_ _05829_ _05832_ _05691_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a22o_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28288_ registers\[2\]\[23\] _10353_ _12528_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18041_ _04808_ _04811_ _04611_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__o21ba_2
XFILLER_173_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_138_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_138_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27239_ _11811_ registers\[37\]\[39\] _11969_ VGND VGND VPWR VPWR _11979_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30250_ registers\[15\]\[26\] _12989_ _13588_ VGND VGND VPWR VPWR _13595_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30181_ _13558_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19992_ registers\[48\]\[46\] registers\[49\]\[46\] registers\[50\]\[46\] registers\[51\]\[46\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__mux4_1
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18943_ registers\[0\]\[16\] registers\[1\]\[16\] registers\[2\]\[16\] registers\[3\]\[16\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux4_1
XFILLER_234_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1410 _00179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1421 _04463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1432 _05039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33940_ clknet_leaf_120_CLK _02054_ VGND VGND VPWR VPWR registers\[37\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_310_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_310_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1443 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18874_ _05618_ _05622_ _05483_ _05484_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o211a_2
XTAP_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1454 _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1465 _05162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17825_ _04602_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_1476 _05485_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33871_ clknet_leaf_133_CLK _01985_ VGND VGND VPWR VPWR registers\[38\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1487 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1498 _07328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35610_ clknet_leaf_15_CLK _03724_ VGND VGND VPWR VPWR registers\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_32822_ clknet_leaf_326_CLK _00936_ VGND VGND VPWR VPWR registers\[55\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_17756_ _04333_ _04533_ _04534_ _04338_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__a22o_1
XFILLER_82_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16707_ registers\[48\]\[18\] registers\[49\]\[18\] registers\[50\]\[18\] registers\[51\]\[18\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15203_ sky130_fd_sc_hd__mux4_1
XFILLER_235_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35541_ clknet_leaf_78_CLK _03655_ VGND VGND VPWR VPWR registers\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_32753_ clknet_leaf_367_CLK _00867_ VGND VGND VPWR VPWR registers\[56\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17687_ registers\[44\]\[46\] registers\[45\]\[46\] registers\[46\]\[46\] registers\[47\]\[46\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__mux4_1
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31704_ _14360_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__clkbuf_1
X_19426_ registers\[36\]\[30\] registers\[37\]\[30\] registers\[38\]\[30\] registers\[39\]\[30\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux4_1
X_35472_ clknet_leaf_137_CLK _03586_ VGND VGND VPWR VPWR registers\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16638_ registers\[52\]\[16\] registers\[53\]\[16\] registers\[54\]\[16\] registers\[55\]\[16\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15136_ sky130_fd_sc_hd__mux4_1
X_32684_ clknet_leaf_371_CLK _00798_ VGND VGND VPWR VPWR registers\[57\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34423_ clknet_leaf_426_CLK _02537_ VGND VGND VPWR VPWR registers\[30\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_31635_ registers\[63\]\[42\] net37 _14321_ VGND VGND VPWR VPWR _14324_ sky130_fd_sc_hd__mux2_1
X_19357_ registers\[56\]\[28\] registers\[57\]\[28\] registers\[58\]\[28\] registers\[59\]\[28\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_377_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_377_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16569_ _14855_ _15067_ _15068_ _14861_ VGND VGND VPWR VPWR _15069_ sky130_fd_sc_hd__a22o_1
X_18308_ registers\[36\]\[0\] registers\[37\]\[0\] registers\[38\]\[0\] registers\[39\]\[0\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__mux4_1
XFILLER_206_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34354_ clknet_leaf_412_CLK _02468_ VGND VGND VPWR VPWR registers\[31\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_31566_ _14287_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__clkbuf_1
X_19288_ registers\[60\]\[26\] registers\[61\]\[26\] registers\[62\]\[26\] registers\[63\]\[26\]
+ _05962_ _05756_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__mux4_1
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33305_ clknet_leaf_29_CLK _01419_ VGND VGND VPWR VPWR registers\[47\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18239_ registers\[28\]\[62\] registers\[29\]\[62\] registers\[30\]\[62\] registers\[31\]\[62\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__mux4_1
X_30517_ _09740_ registers\[13\]\[24\] _13731_ VGND VGND VPWR VPWR _13736_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_129_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_129_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_198_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34285_ clknet_leaf_322_CLK _02399_ VGND VGND VPWR VPWR registers\[32\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_31497_ _14251_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33236_ clknet_leaf_70_CLK _01350_ VGND VGND VPWR VPWR registers\[48\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_36024_ clknet_leaf_332_CLK _04138_ VGND VGND VPWR VPWR registers\[63\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_21250_ _07929_ _07930_ _07931_ _07932_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__a22o_1
X_30448_ _13699_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20201_ _05076_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__clkbuf_8
X_33167_ clknet_leaf_139_CLK _01281_ VGND VGND VPWR VPWR registers\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21181_ _07862_ _07865_ _07730_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__o21ba_2
XFILLER_104_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30379_ _13663_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20132_ registers\[36\]\[50\] registers\[37\]\[50\] registers\[38\]\[50\] registers\[39\]\[50\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__mux4_1
XFILLER_131_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32118_ clknet_leaf_466_CLK _00034_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33098_ clknet_leaf_164_CLK _01212_ VGND VGND VPWR VPWR registers\[51\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20063_ registers\[56\]\[48\] registers\[57\]\[48\] registers\[58\]\[48\] registers\[59\]\[48\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux4_1
X_32049_ clknet_leaf_371_CLK _00227_ VGND VGND VPWR VPWR registers\[62\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_24940_ _09598_ registers\[53\]\[40\] _10702_ VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__mux2_1
XFILLER_225_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_301_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_301_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24871_ _10666_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__clkbuf_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_245_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26610_ _10789_ registers\[41\]\[28\] _11608_ VGND VGND VPWR VPWR _11617_ sky130_fd_sc_hd__mux2_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23822_ _09634_ registers\[29\]\[57\] _10072_ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__mux2_1
XFILLER_2_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35808_ clknet_leaf_484_CLK _03922_ VGND VGND VPWR VPWR registers\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27590_ registers\[34\]\[12\] _10330_ _12162_ VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__mux2_1
XFILLER_85_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26541_ _10856_ registers\[42\]\[60\] _11513_ VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__mux2_1
XANTENNA_318 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20965_ registers\[0\]\[8\] registers\[1\]\[8\] registers\[2\]\[8\] registers\[3\]\[8\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__mux4_1
X_35739_ clknet_leaf_480_CLK _03853_ VGND VGND VPWR VPWR registers\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_23753_ _09565_ registers\[29\]\[24\] _10039_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__mux2_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _07372_ _09343_ _09344_ _07382_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__a22o_1
X_29260_ _13074_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26472_ _10787_ registers\[42\]\[27\] _11536_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23684_ registers\[61\]\[57\] _09813_ _09998_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__mux2_1
X_20896_ _07366_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__buf_4
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28211_ _12491_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__clkbuf_1
X_25423_ _10827_ registers\[50\]\[46\] _10981_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__mux2_1
X_22635_ registers\[40\]\[56\] registers\[41\]\[56\] registers\[42\]\[56\] registers\[43\]\[56\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__mux4_1
X_29191_ net40 VGND VGND VPWR VPWR _13029_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_368_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_368_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28142_ _11767_ registers\[30\]\[18\] _12446_ VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__mux2_1
X_22566_ registers\[20\]\[53\] registers\[21\]\[53\] registers\[22\]\[53\] registers\[23\]\[53\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__mux4_1
X_25354_ _10758_ registers\[50\]\[13\] _10948_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__mux2_1
XFILLER_166_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_934 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24305_ registers\[57\]\[19\] _10344_ _10326_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__mux2_1
X_21517_ _08126_ _08190_ _08191_ _08129_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__a22o_1
X_28073_ _12418_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_1
X_22497_ _09109_ _09143_ _09144_ _09114_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__a22o_1
X_25285_ _10825_ registers\[51\]\[45\] _10909_ VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__mux2_1
XFILLER_181_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27024_ _11866_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_1
X_24236_ _09640_ registers\[58\]\[60\] _10232_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__mux2_1
X_21448_ _08119_ _08122_ _08123_ _08124_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__a22o_1
XFILLER_182_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24167_ _09571_ registers\[58\]\[27\] _10255_ VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__mux2_1
X_21379_ _07983_ _08056_ _08057_ _07989_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__a22o_1
XFILLER_162_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23118_ _09657_ VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__clkbuf_8
X_24098_ _09638_ registers\[5\]\[59\] _10216_ VGND VGND VPWR VPWR _10226_ sky130_fd_sc_hd__mux2_1
XFILLER_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28975_ registers\[24\]\[29\] _10365_ _12883_ VGND VGND VPWR VPWR _12893_ sky130_fd_sc_hd__mux2_1
X_23049_ _09629_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27926_ _12341_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27857_ _12305_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ registers\[16\]\[43\] registers\[17\]\[43\] registers\[18\]\[43\] registers\[19\]\[43\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__mux4_1
X_26808_ _11721_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__clkbuf_1
XTAP_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ registers\[0\]\[6\] registers\[1\]\[6\] registers\[2\]\[6\] registers\[3\]\[6\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__mux4_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27788_ registers\[33\]\[42\] _10393_ _12266_ VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__mux2_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29527_ registers\[20\]\[3\] _12941_ _13211_ VGND VGND VPWR VPWR _13215_ sky130_fd_sc_hd__mux2_1
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _04289_ _04325_ _04326_ _04292_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__a22o_1
XFILLER_217_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26739_ _11685_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_830 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_841 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_852 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29458_ _13178_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17472_ _15946_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_863 _09335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_874 _09523_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19211_ _05950_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16423_ _14920_ _14925_ _14926_ VGND VGND VPWR VPWR _14927_ sky130_fd_sc_hd__o21ba_1
XANTENNA_885 _09588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28409_ _12595_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_896 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29389_ _13142_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_359_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_359_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31420_ _09666_ registers\[6\]\[4\] _14206_ VGND VGND VPWR VPWR _14211_ sky130_fd_sc_hd__mux2_1
X_19142_ _05076_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__clkbuf_4
XFILLER_242_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16354_ registers\[48\]\[8\] registers\[49\]\[8\] registers\[50\]\[8\] registers\[51\]\[8\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _14860_ sky130_fd_sc_hd__mux4_1
XFILLER_157_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31351_ _14174_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__clkbuf_1
X_19073_ registers\[36\]\[20\] registers\[37\]\[20\] registers\[38\]\[20\] registers\[39\]\[20\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__mux4_1
XFILLER_146_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16285_ registers\[52\]\[6\] registers\[53\]\[6\] registers\[54\]\[6\] registers\[55\]\[6\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14793_ sky130_fd_sc_hd__mux4_1
XFILLER_201_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30302_ _13622_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__clkbuf_1
X_18024_ _04486_ _04794_ _04795_ _04489_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a22o_1
X_34070_ clknet_leaf_120_CLK _02184_ VGND VGND VPWR VPWR registers\[35\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31282_ _14138_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__clkbuf_1
X_33021_ clknet_leaf_290_CLK _01135_ VGND VGND VPWR VPWR registers\[52\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_30233_ registers\[15\]\[18\] _12972_ _13577_ VGND VGND VPWR VPWR _13586_ sky130_fd_sc_hd__mux2_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30164_ _13549_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19975_ registers\[24\]\[45\] registers\[25\]\[45\] registers\[26\]\[45\] registers\[27\]\[45\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__mux4_1
XFILLER_80_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18926_ registers\[32\]\[16\] registers\[33\]\[16\] registers\[34\]\[16\] registers\[35\]\[16\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__mux4_1
XFILLER_136_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34972_ clknet_leaf_492_CLK _03086_ VGND VGND VPWR VPWR registers\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_30095_ _13513_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1240 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1251 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1262 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33923_ clknet_leaf_254_CLK _02037_ VGND VGND VPWR VPWR registers\[38\]\[53\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1273 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1284 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18857_ _05583_ _05590_ _05599_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or4_2
XFILLER_80_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1295 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17808_ _04548_ _04584_ _04585_ _04552_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a22o_1
XFILLER_212_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33854_ clknet_leaf_296_CLK _01968_ VGND VGND VPWR VPWR registers\[3\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_18788_ _05539_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17739_ registers\[0\]\[47\] registers\[1\]\[47\] registers\[2\]\[47\] registers\[3\]\[47\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__mux4_1
X_32805_ clknet_leaf_442_CLK _00919_ VGND VGND VPWR VPWR registers\[55\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30997_ registers\[10\]\[60\] _13060_ _13921_ VGND VGND VPWR VPWR _13988_ sky130_fd_sc_hd__mux2_1
X_33785_ clknet_leaf_338_CLK _01899_ VGND VGND VPWR VPWR registers\[40\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35524_ clknet_6_60__leaf_CLK _03638_ VGND VGND VPWR VPWR registers\[13\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_20750_ registers\[48\]\[2\] registers\[49\]\[2\] registers\[50\]\[2\] registers\[51\]\[2\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32736_ clknet_leaf_44_CLK _00850_ VGND VGND VPWR VPWR registers\[56\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19409_ _06036_ _06141_ _06142_ _06039_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__a22o_1
X_20681_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__buf_4
X_35455_ clknet_leaf_197_CLK _03569_ VGND VGND VPWR VPWR registers\[14\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_32667_ clknet_leaf_35_CLK _00781_ VGND VGND VPWR VPWR registers\[57\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22420_ registers\[28\]\[49\] registers\[29\]\[49\] registers\[30\]\[49\] registers\[31\]\[49\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__mux4_1
XFILLER_17_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31618_ registers\[63\]\[34\] net28 _14310_ VGND VGND VPWR VPWR _14315_ sky130_fd_sc_hd__mux2_1
X_34406_ clknet_leaf_448_CLK _02520_ VGND VGND VPWR VPWR registers\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32598_ clknet_leaf_65_CLK _00712_ VGND VGND VPWR VPWR registers\[58\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35386_ clknet_leaf_302_CLK _03500_ VGND VGND VPWR VPWR registers\[15\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22351_ _08999_ _09002_ _08773_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__o21ba_1
X_31549_ registers\[63\]\[1\] net12 _14277_ VGND VGND VPWR VPWR _14279_ sky130_fd_sc_hd__mux2_1
XFILLER_137_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34337_ clknet_leaf_488_CLK _02451_ VGND VGND VPWR VPWR registers\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_21302_ _07312_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__clkbuf_4
X_25070_ _10783_ registers\[52\]\[25\] _10773_ VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__mux2_1
X_22282_ _08912_ _08919_ _08928_ _08935_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__or4_4
X_34268_ clknet_leaf_23_CLK _02382_ VGND VGND VPWR VPWR registers\[32\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24021_ _09561_ registers\[5\]\[22\] _10183_ VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33219_ clknet_leaf_232_CLK _01333_ VGND VGND VPWR VPWR registers\[4\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_36007_ clknet_leaf_437_CLK _04121_ VGND VGND VPWR VPWR registers\[63\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21233_ registers\[48\]\[16\] registers\[49\]\[16\] registers\[50\]\[16\] registers\[51\]\[16\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__mux4_1
X_34199_ clknet_leaf_109_CLK _02313_ VGND VGND VPWR VPWR registers\[33\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_942 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21164_ _07783_ _07847_ _07848_ _07786_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__a22o_1
XFILLER_131_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ _06722_ _06827_ _06828_ _06725_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__a22o_1
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28760_ _11845_ registers\[26\]\[55\] _12774_ VGND VGND VPWR VPWR _12780_ sky130_fd_sc_hd__mux2_1
X_25972_ _10827_ registers\[46\]\[46\] _11274_ VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__mux2_1
X_21095_ _07776_ _07779_ _07780_ _07781_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__a22o_1
XFILLER_154_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27711_ _12228_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_1
X_20046_ registers\[16\]\[47\] registers\[17\]\[47\] registers\[18\]\[47\] registers\[19\]\[47\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__mux4_1
X_24923_ _09582_ registers\[53\]\[32\] _10691_ VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__mux2_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28691_ _11776_ registers\[26\]\[22\] _12741_ VGND VGND VPWR VPWR _12744_ sky130_fd_sc_hd__mux2_1
XFILLER_218_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27642_ registers\[34\]\[37\] _10382_ _12184_ VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__mux2_1
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24854_ _10015_ _10512_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__nand2_8
XFILLER_74_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _09617_ registers\[29\]\[49\] _10061_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__mux2_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27573_ registers\[34\]\[4\] _10313_ _12151_ VGND VGND VPWR VPWR _12156_ sky130_fd_sc_hd__mux2_1
XANTENNA_104 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24785_ _10621_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _08423_ _08657_ _08658_ _08428_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__a22o_1
XANTENNA_137 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29312_ _13101_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26524_ _11571_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _09548_ registers\[29\]\[16\] _10028_ VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__mux2_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20948_ _07635_ _07638_ _07310_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__o21ba_2
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_159 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29243_ net59 VGND VGND VPWR VPWR _13064_ sky130_fd_sc_hd__buf_2
XFILLER_144_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26455_ _10770_ registers\[42\]\[19\] _11525_ VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__mux2_1
XFILLER_202_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23667_ registers\[61\]\[49\] _09795_ _09987_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__mux2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20879_ registers\[56\]\[6\] registers\[57\]\[6\] registers\[58\]\[6\] registers\[59\]\[6\]
+ _07508_ _07317_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__mux4_1
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25406_ _10810_ registers\[50\]\[38\] _10970_ VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__mux2_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22618_ _09258_ _09261_ _09091_ _09092_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__o211a_1
X_29174_ _13017_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26386_ _10835_ registers\[43\]\[50\] _11498_ VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__mux2_1
XFILLER_201_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23598_ registers\[61\]\[16\] _09691_ _09954_ VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__mux2_1
X_28125_ _12434_ VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__buf_4
XFILLER_220_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25337_ _10741_ registers\[50\]\[5\] _10937_ VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__mux2_1
X_22549_ registers\[60\]\[53\] registers\[61\]\[53\] registers\[62\]\[53\] registers\[63\]\[53\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__mux4_1
XFILLER_220_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16070_ net69 net70 VGND VGND VPWR VPWR _14584_ sky130_fd_sc_hd__or2_4
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28056_ _11816_ registers\[31\]\[41\] _12408_ VGND VGND VPWR VPWR _12410_ sky130_fd_sc_hd__mux2_1
X_25268_ _10808_ registers\[51\]\[37\] _10898_ VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__mux2_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27007_ _11854_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24219_ _10290_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25199_ _10739_ registers\[51\]\[4\] _10865_ VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__mux2_1
XFILLER_151_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16972_ registers\[28\]\[25\] registers\[29\]\[25\] registers\[30\]\[25\] registers\[31\]\[25\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15461_ sky130_fd_sc_hd__mux4_1
X_19760_ registers\[12\]\[39\] registers\[13\]\[39\] registers\[14\]\[39\] registers\[15\]\[39\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__mux4_1
XFILLER_150_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28958_ _12884_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18711_ _05461_ _05464_ _05163_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__o21ba_1
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19691_ _06413_ _06416_ _06180_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__o21ba_1
X_27909_ _12332_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__clkbuf_1
X_28889_ _11839_ registers\[25\]\[52\] _12845_ VGND VGND VPWR VPWR _12848_ sky130_fd_sc_hd__mux2_1
XFILLER_232_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18642_ registers\[40\]\[8\] registers\[41\]\[8\] registers\[42\]\[8\] registers\[43\]\[8\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__mux4_1
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30920_ registers\[10\]\[23\] _12983_ _13944_ VGND VGND VPWR VPWR _13948_ sky130_fd_sc_hd__mux2_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30851_ _13911_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__clkbuf_1
X_18573_ registers\[32\]\[6\] registers\[33\]\[6\] registers\[34\]\[6\] registers\[35\]\[6\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__mux4_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17524_ _04306_ _04309_ _15955_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__o21ba_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33570_ clknet_leaf_56_CLK _01684_ VGND VGND VPWR VPWR registers\[43\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_233_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30782_ _13875_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_660 _05297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32521_ clknet_leaf_162_CLK _00635_ VGND VGND VPWR VPWR registers\[60\]\[59\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_671 _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_682 _06152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17455_ _15892_ _15928_ _15929_ _15896_ VGND VGND VPWR VPWR _15930_ sky130_fd_sc_hd__a22o_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_693 _06919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16406_ registers\[16\]\[9\] registers\[17\]\[9\] registers\[18\]\[9\] registers\[19\]\[9\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14911_ sky130_fd_sc_hd__mux4_1
X_32452_ clknet_leaf_203_CLK _00566_ VGND VGND VPWR VPWR registers\[29\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_35240_ clknet_leaf_405_CLK _03354_ VGND VGND VPWR VPWR registers\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_17386_ registers\[0\]\[37\] registers\[1\]\[37\] registers\[2\]\[37\] registers\[3\]\[37\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15863_ sky130_fd_sc_hd__mux4_1
X_31403_ _14201_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__clkbuf_1
X_19125_ _05863_ _05866_ _05826_ _05827_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__o211a_1
X_16337_ registers\[20\]\[7\] registers\[21\]\[7\] registers\[22\]\[7\] registers\[23\]\[7\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14844_ sky130_fd_sc_hd__mux4_1
XFILLER_119_928 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35171_ clknet_leaf_474_CLK _03285_ VGND VGND VPWR VPWR registers\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32383_ clknet_leaf_293_CLK _00497_ VGND VGND VPWR VPWR registers\[61\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34122_ clknet_leaf_156_CLK _02236_ VGND VGND VPWR VPWR registers\[35\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19056_ _05693_ _05798_ _05799_ _05696_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__a22o_1
X_31334_ _14165_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__clkbuf_1
X_16268_ _14601_ _14775_ _14776_ _14611_ VGND VGND VPWR VPWR _14777_ sky130_fd_sc_hd__a22o_1
XFILLER_161_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18007_ _04676_ _04777_ _04778_ _04681_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__a22o_1
X_34053_ clknet_leaf_260_CLK _02167_ VGND VGND VPWR VPWR registers\[36\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_31265_ registers\[8\]\[59\] net55 _14119_ VGND VGND VPWR VPWR _14129_ sky130_fd_sc_hd__mux2_1
XFILLER_173_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16199_ _14588_ _14708_ _14709_ _14598_ VGND VGND VPWR VPWR _14710_ sky130_fd_sc_hd__a22o_1
XFILLER_142_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_60_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33004_ clknet_leaf_371_CLK _01118_ VGND VGND VPWR VPWR registers\[52\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30216_ _13565_ VGND VGND VPWR VPWR _13577_ sky130_fd_sc_hd__buf_4
XFILLER_160_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31196_ registers\[8\]\[26\] net19 _14086_ VGND VGND VPWR VPWR _14093_ sky130_fd_sc_hd__mux2_1
XFILLER_102_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30147_ registers\[16\]\[41\] _13021_ _13539_ VGND VGND VPWR VPWR _13541_ sky130_fd_sc_hd__mux2_1
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19958_ _06672_ _06675_ _06504_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18909_ registers\[8\]\[15\] registers\[9\]\[15\] registers\[10\]\[15\] registers\[11\]\[15\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__mux4_1
X_34955_ clknet_leaf_143_CLK _03069_ VGND VGND VPWR VPWR registers\[22\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_30078_ _13504_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1070 _14347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19889_ registers\[44\]\[43\] registers\[45\]\[43\] registers\[46\]\[43\] registers\[47\]\[43\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__mux4_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1081 _14496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1092 _14520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21920_ _08272_ _08582_ _08583_ _08275_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__a22o_1
X_33906_ clknet_leaf_356_CLK _02020_ VGND VGND VPWR VPWR registers\[38\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34886_ clknet_leaf_208_CLK _03000_ VGND VGND VPWR VPWR registers\[23\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_243_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33837_ clknet_leaf_388_CLK _01951_ VGND VGND VPWR VPWR registers\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_21851_ _07305_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__buf_4
XFILLER_83_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20802_ _07386_ _07496_ _07497_ _07396_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__a22o_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24570_ _10505_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21782_ registers\[12\]\[31\] registers\[13\]\[31\] registers\[14\]\[31\] registers\[15\]\[31\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__mux4_1
XFILLER_24_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33768_ clknet_leaf_430_CLK _01882_ VGND VGND VPWR VPWR registers\[40\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23521_ _09919_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__clkbuf_1
X_35507_ clknet_leaf_355_CLK _03621_ VGND VGND VPWR VPWR registers\[13\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20733_ _07427_ _07430_ _07399_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__o21ba_1
X_32719_ clknet_leaf_173_CLK _00833_ VGND VGND VPWR VPWR registers\[56\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33699_ clknet_leaf_55_CLK _01813_ VGND VGND VPWR VPWR registers\[41\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26240_ _10825_ registers\[44\]\[45\] _11416_ VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__mux2_1
X_35438_ clknet_leaf_393_CLK _03552_ VGND VGND VPWR VPWR registers\[14\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_23452_ _09883_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
X_20664_ _07316_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22403_ registers\[56\]\[49\] registers\[57\]\[49\] registers\[58\]\[49\] registers\[59\]\[49\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__mux4_1
XFILLER_137_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23383_ _09845_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
X_26171_ _10756_ registers\[44\]\[12\] _11383_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__mux2_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20595_ _07293_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__buf_2
XFILLER_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35369_ clknet_leaf_398_CLK _03483_ VGND VGND VPWR VPWR registers\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25122_ net37 VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__buf_2
XFILLER_192_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22334_ registers\[60\]\[47\] registers\[61\]\[47\] registers\[62\]\[47\] registers\[63\]\[47\]
+ _08884_ _08678_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__mux4_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29930_ registers\[17\]\[2\] _12939_ _13424_ VGND VGND VPWR VPWR _13427_ sky130_fd_sc_hd__mux2_1
X_22265_ _08915_ _08918_ _08748_ _08749_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__o211a_1
X_25053_ net13 VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_51_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24004_ _09544_ registers\[5\]\[14\] _10172_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__mux2_1
X_21216_ registers\[24\]\[15\] registers\[25\]\[15\] registers\[26\]\[15\] registers\[27\]\[15\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__mux4_1
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29861_ _13390_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__clkbuf_1
X_22196_ registers\[60\]\[43\] registers\[61\]\[43\] registers\[62\]\[43\] registers\[63\]\[43\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__mux4_1
XFILLER_132_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28812_ _12807_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__clkbuf_1
X_21147_ registers\[4\]\[13\] registers\[5\]\[13\] registers\[6\]\[13\] registers\[7\]\[13\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__mux4_1
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29792_ _13354_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28743_ _11828_ registers\[26\]\[47\] _12763_ VGND VGND VPWR VPWR _12771_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21078_ _07586_ _07764_ _07765_ _07589_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__a22o_1
X_25955_ _10810_ registers\[46\]\[38\] _11263_ VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__mux2_1
XFILLER_246_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20029_ _06576_ _06741_ _06744_ _06579_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__a22o_1
XFILLER_4_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24906_ _09565_ registers\[53\]\[24\] _10680_ VGND VGND VPWR VPWR _10685_ sky130_fd_sc_hd__mux2_1
XFILLER_207_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28674_ _11759_ registers\[26\]\[14\] _12730_ VGND VGND VPWR VPWR _12735_ sky130_fd_sc_hd__mux2_1
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25886_ _10741_ registers\[46\]\[5\] _11230_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__mux2_1
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27625_ registers\[34\]\[29\] _10365_ _12173_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__mux2_1
XFILLER_98_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24837_ _10648_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27556_ _12145_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24768_ _10612_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26507_ _11562_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__clkbuf_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23719_ _09531_ registers\[29\]\[8\] _10017_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__mux2_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27487_ _12109_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24699_ _09630_ registers\[55\]\[55\] _10569_ VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__mux2_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29226_ registers\[23\]\[56\] _13052_ _13040_ VGND VGND VPWR VPWR _13053_ sky130_fd_sc_hd__mux2_1
X_17240_ registers\[56\]\[33\] registers\[57\]\[33\] registers\[58\]\[33\] registers\[59\]\[33\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15721_ sky130_fd_sc_hd__mux4_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26438_ _11526_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__clkbuf_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29157_ net28 VGND VGND VPWR VPWR _13006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17171_ _15650_ _15653_ _15612_ VGND VGND VPWR VPWR _15654_ sky130_fd_sc_hd__o21ba_1
X_26369_ _10819_ registers\[43\]\[42\] _11487_ VGND VGND VPWR VPWR _11490_ sky130_fd_sc_hd__mux2_1
X_16122_ _14558_ _14633_ _14634_ _14568_ VGND VGND VPWR VPWR _14635_ sky130_fd_sc_hd__a22o_1
X_28108_ _12437_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__clkbuf_1
X_29088_ _12959_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16053_ _14499_ VGND VGND VPWR VPWR _14567_ sky130_fd_sc_hd__buf_12
XFILLER_109_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28039_ _11799_ registers\[31\]\[33\] _12397_ VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_42_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_48__f_CLK clknet_5_24_0_CLK VGND VGND VPWR VPWR clknet_6_48__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31050_ _14016_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30001_ registers\[17\]\[36\] _13010_ _13457_ VGND VGND VPWR VPWR _13464_ sky130_fd_sc_hd__mux2_1
X_19812_ _05130_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_116_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19743_ _05069_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__buf_4
XFILLER_172_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16955_ _15198_ _15442_ _15443_ _15204_ VGND VGND VPWR VPWR _15444_ sky130_fd_sc_hd__a22o_1
XFILLER_133_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34740_ clknet_leaf_413_CLK _02854_ VGND VGND VPWR VPWR registers\[25\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31952_ clknet_leaf_492_CLK _00150_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
X_16886_ _15373_ _15376_ _15269_ VGND VGND VPWR VPWR _15377_ sky130_fd_sc_hd__o21ba_1
X_19674_ _05122_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18625_ _05377_ _05380_ _05103_ _05105_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__o211a_1
X_30903_ registers\[10\]\[15\] _12966_ _13933_ VGND VGND VPWR VPWR _13939_ sky130_fd_sc_hd__mux2_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31883_ _14454_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__clkbuf_1
X_34671_ clknet_leaf_410_CLK _02785_ VGND VGND VPWR VPWR registers\[26\]\[33\] sky130_fd_sc_hd__dfxtp_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33622_ clknet_leaf_126_CLK _01736_ VGND VGND VPWR VPWR registers\[42\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_30834_ _13902_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18556_ registers\[8\]\[5\] registers\[9\]\[5\] registers\[10\]\[5\] registers\[11\]\[5\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__mux4_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17507_ _14510_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__clkbuf_4
X_33553_ clknet_leaf_129_CLK _01667_ VGND VGND VPWR VPWR registers\[43\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_18487_ _05243_ _05246_ _05103_ _05105_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__o211a_1
X_30765_ _13866_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_490 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32504_ clknet_leaf_332_CLK _00618_ VGND VGND VPWR VPWR registers\[60\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17438_ _15910_ _15913_ _15645_ VGND VGND VPWR VPWR _15914_ sky130_fd_sc_hd__o21ba_1
X_33484_ clknet_leaf_164_CLK _01598_ VGND VGND VPWR VPWR registers\[45\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30696_ registers\[12\]\[45\] _13029_ _13824_ VGND VGND VPWR VPWR _13830_ sky130_fd_sc_hd__mux2_1
XANTENNA_15 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35223_ clknet_leaf_92_CLK _03337_ VGND VGND VPWR VPWR registers\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_32435_ clknet_leaf_412_CLK _00549_ VGND VGND VPWR VPWR registers\[29\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_17369_ registers\[40\]\[37\] registers\[41\]\[37\] registers\[42\]\[37\] registers\[43\]\[37\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15846_ sky130_fd_sc_hd__mux4_1
XFILLER_203_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19108_ _05162_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__buf_2
X_20380_ registers\[0\]\[57\] registers\[1\]\[57\] registers\[2\]\[57\] registers\[3\]\[57\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__mux4_1
XFILLER_192_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35154_ clknet_leaf_101_CLK _03268_ VGND VGND VPWR VPWR registers\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_32366_ clknet_leaf_370_CLK _00480_ VGND VGND VPWR VPWR registers\[61\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34105_ clknet_leaf_337_CLK _02219_ VGND VGND VPWR VPWR registers\[35\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31317_ _14156_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__clkbuf_1
X_19039_ _05540_ _05779_ _05782_ _05545_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__a22o_1
X_35085_ clknet_leaf_145_CLK _03199_ VGND VGND VPWR VPWR registers\[20\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32297_ clknet_leaf_408_CLK _00411_ VGND VGND VPWR VPWR registers\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xoutput100 net100 VGND VGND VPWR VPWR D1[19] sky130_fd_sc_hd__buf_2
Xoutput111 net111 VGND VGND VPWR VPWR D1[29] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_33_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_33_CLK sky130_fd_sc_hd__clkbuf_16
Xoutput122 net122 VGND VGND VPWR VPWR D1[39] sky130_fd_sc_hd__buf_2
X_22050_ registers\[56\]\[39\] registers\[57\]\[39\] registers\[58\]\[39\] registers\[59\]\[39\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__mux4_1
Xoutput133 net133 VGND VGND VPWR VPWR D1[49] sky130_fd_sc_hd__buf_2
X_31248_ _14120_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34036_ clknet_leaf_344_CLK _02150_ VGND VGND VPWR VPWR registers\[36\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput144 net144 VGND VGND VPWR VPWR D1[59] sky130_fd_sc_hd__buf_2
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput155 net155 VGND VGND VPWR VPWR D2[10] sky130_fd_sc_hd__buf_2
XFILLER_216_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput166 net166 VGND VGND VPWR VPWR D2[20] sky130_fd_sc_hd__buf_2
X_21001_ registers\[12\]\[9\] registers\[13\]\[9\] registers\[14\]\[9\] registers\[15\]\[9\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__mux4_1
XFILLER_99_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 net177 VGND VGND VPWR VPWR D2[30] sky130_fd_sc_hd__buf_2
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput188 net188 VGND VGND VPWR VPWR D2[40] sky130_fd_sc_hd__buf_2
XFILLER_87_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31179_ registers\[8\]\[18\] net10 _14075_ VGND VGND VPWR VPWR _14084_ sky130_fd_sc_hd__mux2_1
Xoutput199 net199 VGND VGND VPWR VPWR D2[50] sky130_fd_sc_hd__buf_2
XFILLER_153_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35987_ clknet_leaf_182_CLK _04101_ VGND VGND VPWR VPWR registers\[63\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25740_ _11158_ VGND VGND VPWR VPWR _11159_ sky130_fd_sc_hd__buf_4
XFILLER_96_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34938_ clknet_leaf_308_CLK _03052_ VGND VGND VPWR VPWR registers\[22\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22952_ _09563_ registers\[62\]\[23\] _09557_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__mux2_1
XFILLER_110_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21903_ registers\[36\]\[35\] registers\[37\]\[35\] registers\[38\]\[35\] registers\[39\]\[35\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__mux4_1
X_25671_ registers\[48\]\[32\] _10372_ _11119_ VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__mux2_1
X_22883_ net12 VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__clkbuf_4
X_34869_ clknet_leaf_386_CLK _02983_ VGND VGND VPWR VPWR registers\[23\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27410_ registers\[36\]\[56\] _10422_ _12062_ VGND VGND VPWR VPWR _12069_ sky130_fd_sc_hd__mux2_1
X_24622_ _10534_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
X_28390_ _12585_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21834_ registers\[32\]\[33\] registers\[33\]\[33\] registers\[34\]\[33\] registers\[35\]\[33\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__mux4_1
XFILLER_110_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27341_ registers\[36\]\[23\] _10353_ _12029_ VGND VGND VPWR VPWR _12033_ sky130_fd_sc_hd__mux2_1
X_24553_ _09622_ registers\[56\]\[51\] _10495_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__mux2_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21765_ registers\[40\]\[31\] registers\[41\]\[31\] registers\[42\]\[31\] registers\[43\]\[31\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__mux4_1
XFILLER_197_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23504_ _09910_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__clkbuf_1
X_27272_ _11996_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20716_ registers\[60\]\[1\] registers\[61\]\[1\] registers\[62\]\[1\] registers\[63\]\[1\]
+ _07327_ _07329_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__mux4_1
XFILLER_145_1267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24484_ _10460_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
X_21696_ _08362_ _08365_ _08054_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__o21ba_1
X_29011_ registers\[24\]\[46\] _10401_ _12905_ VGND VGND VPWR VPWR _12912_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26223_ _10808_ registers\[44\]\[37\] _11405_ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__mux2_1
X_23435_ _09874_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
X_20647_ registers\[8\]\[0\] registers\[9\]\[0\] registers\[10\]\[0\] registers\[11\]\[0\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__mux4_1
XFILLER_109_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26154_ _10739_ registers\[44\]\[4\] _11372_ VGND VGND VPWR VPWR _11377_ sky130_fd_sc_hd__mux2_1
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20578_ net71 VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__buf_6
XFILLER_221_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23366_ _09836_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_3_0_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_3_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25105_ _10807_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__clkbuf_1
X_22317_ registers\[20\]\[46\] registers\[21\]\[46\] registers\[22\]\[46\] registers\[23\]\[46\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__mux4_1
XFILLER_139_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26085_ _11340_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
X_23297_ net43 VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__clkbuf_4
XFILLER_139_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_24_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29913_ _13417_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25036_ _10760_ registers\[52\]\[14\] _10752_ VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__mux2_1
XFILLER_191_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22248_ _08766_ _08901_ _08902_ _08771_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__a22o_1
XFILLER_180_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22179_ _07363_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__buf_4
X_29844_ _13381_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29775_ registers\[1\]\[57\] _13054_ _13337_ VGND VGND VPWR VPWR _13345_ sky130_fd_sc_hd__mux2_1
X_26987_ net49 VGND VGND VPWR VPWR _11841_ sky130_fd_sc_hd__buf_4
XFILLER_28_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16740_ registers\[44\]\[19\] registers\[45\]\[19\] registers\[46\]\[19\] registers\[47\]\[19\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15235_ sky130_fd_sc_hd__mux4_1
XFILLER_115_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28726_ _11811_ registers\[26\]\[39\] _12752_ VGND VGND VPWR VPWR _12762_ sky130_fd_sc_hd__mux2_1
X_25938_ _11229_ VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__buf_4
XFILLER_247_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28657_ _11742_ registers\[26\]\[6\] _12719_ VGND VGND VPWR VPWR _12726_ sky130_fd_sc_hd__mux2_1
X_16671_ _15162_ _15167_ _14926_ VGND VGND VPWR VPWR _15168_ sky130_fd_sc_hd__o21ba_1
X_25869_ _11226_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18410_ registers\[36\]\[1\] registers\[37\]\[1\] registers\[38\]\[1\] registers\[39\]\[1\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux4_1
XFILLER_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19390_ _05069_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__buf_4
X_27608_ _12174_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28588_ _12689_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__clkbuf_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18341_ net82 VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__buf_12
XFILLER_167_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27539_ _11841_ registers\[35\]\[53\] _12133_ VGND VGND VPWR VPWR _12137_ sky130_fd_sc_hd__mux2_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _05032_ _05035_ _14613_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__o21ba_1
XFILLER_187_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30550_ _13708_ VGND VGND VPWR VPWR _13753_ sky130_fd_sc_hd__buf_4
XFILLER_202_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17223_ registers\[16\]\[32\] registers\[17\]\[32\] registers\[18\]\[32\] registers\[19\]\[32\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15705_ sky130_fd_sc_hd__mux4_1
XFILLER_198_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29209_ _13041_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30481_ _09672_ registers\[13\]\[7\] _13709_ VGND VGND VPWR VPWR _13717_ sky130_fd_sc_hd__mux2_1
XFILLER_156_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 DW[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_6
X_32220_ clknet_leaf_237_CLK _00334_ VGND VGND VPWR VPWR registers\[9\]\[51\] sky130_fd_sc_hd__dfxtp_1
Xinput24 DW[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
X_17154_ _14600_ VGND VGND VPWR VPWR _15638_ sky130_fd_sc_hd__clkbuf_4
Xinput35 DW[40] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
Xinput46 DW[50] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_6
Xinput57 DW[60] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_16
Xinput68 R1[3] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_8
X_16105_ registers\[32\]\[1\] registers\[33\]\[1\] registers\[34\]\[1\] registers\[35\]\[1\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14618_ sky130_fd_sc_hd__mux4_1
XFILLER_128_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32151_ clknet_leaf_117_CLK _00265_ VGND VGND VPWR VPWR registers\[39\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xinput79 R3[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
X_17085_ _15567_ _15570_ _15302_ VGND VGND VPWR VPWR _15571_ sky130_fd_sc_hd__o21ba_1
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_15_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31102_ _14043_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__clkbuf_1
X_16036_ registers\[52\]\[0\] registers\[53\]\[0\] registers\[54\]\[0\] registers\[55\]\[0\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14550_ sky130_fd_sc_hd__mux4_1
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32082_ clknet_leaf_490_CLK _00044_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35910_ clknet_leaf_210_CLK _04024_ VGND VGND VPWR VPWR registers\[7\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_31033_ _14007_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35841_ clknet_leaf_237_CLK _03955_ VGND VGND VPWR VPWR registers\[8\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_17987_ registers\[8\]\[54\] registers\[9\]\[54\] registers\[10\]\[54\] registers\[11\]\[54\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux4_1
XFILLER_211_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19726_ registers\[12\]\[38\] registers\[13\]\[38\] registers\[14\]\[38\] registers\[15\]\[38\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__mux4_1
X_35772_ clknet_leaf_301_CLK _03886_ VGND VGND VPWR VPWR registers\[0\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16938_ registers\[16\]\[24\] registers\[17\]\[24\] registers\[18\]\[24\] registers\[19\]\[24\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15428_ sky130_fd_sc_hd__mux4_1
X_32984_ clknet_leaf_53_CLK _01098_ VGND VGND VPWR VPWR registers\[52\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34723_ clknet_leaf_445_CLK _02837_ VGND VGND VPWR VPWR registers\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_31935_ _14481_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__clkbuf_1
X_19657_ _06378_ _06383_ _06180_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__o21ba_1
XFILLER_77_1106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16869_ registers\[24\]\[22\] registers\[25\]\[22\] registers\[26\]\[22\] registers\[27\]\[22\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15361_ sky130_fd_sc_hd__mux4_1
XFILLER_52_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18608_ _05335_ _05344_ _05355_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or4_4
X_34654_ clknet_leaf_4_CLK _02768_ VGND VGND VPWR VPWR registers\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19588_ _05111_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__buf_6
X_31866_ _14445_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33605_ clknet_leaf_250_CLK _01719_ VGND VGND VPWR VPWR registers\[43\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18539_ _05297_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__clkbuf_1
X_30817_ _13893_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__clkbuf_1
X_31797_ registers\[59\]\[55\] net51 _14403_ VGND VGND VPWR VPWR _14409_ sky130_fd_sc_hd__mux2_1
X_34585_ clknet_leaf_21_CLK _02699_ VGND VGND VPWR VPWR registers\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33536_ clknet_leaf_257_CLK _01650_ VGND VGND VPWR VPWR registers\[44\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_21550_ registers\[36\]\[25\] registers\[37\]\[25\] registers\[38\]\[25\] registers\[39\]\[25\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__mux4_1
X_30748_ _13857_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20501_ _05040_ _07201_ _07202_ _05050_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__a22o_1
X_21481_ registers\[32\]\[23\] registers\[33\]\[23\] registers\[34\]\[23\] registers\[35\]\[23\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__mux4_1
X_33467_ clknet_leaf_278_CLK _01581_ VGND VGND VPWR VPWR registers\[45\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_30679_ registers\[12\]\[37\] _13012_ _13813_ VGND VGND VPWR VPWR _13821_ sky130_fd_sc_hd__mux2_1
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35206_ clknet_leaf_153_CLK _03320_ VGND VGND VPWR VPWR registers\[18\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20432_ registers\[56\]\[59\] registers\[57\]\[59\] registers\[58\]\[59\] registers\[59\]\[59\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__mux4_1
X_23220_ net18 VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32418_ clknet_leaf_473_CLK _00532_ VGND VGND VPWR VPWR registers\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_36186_ clknet_leaf_92_CLK _00067_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33398_ clknet_leaf_340_CLK _01512_ VGND VGND VPWR VPWR registers\[46\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35137_ clknet_leaf_240_CLK _03251_ VGND VGND VPWR VPWR registers\[1\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_20363_ _07048_ _07055_ _07062_ _07069_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__or4_2
XFILLER_179_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23151_ _09701_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32349_ clknet_leaf_55_CLK _00463_ VGND VGND VPWR VPWR registers\[61\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22102_ _07275_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__clkbuf_4
XTAP_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23082_ _09652_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__buf_8
X_20294_ _05111_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__buf_6
XFILLER_162_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35068_ clknet_leaf_307_CLK _03182_ VGND VGND VPWR VPWR registers\[20\]\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_6_31__f_CLK clknet_5_15_0_CLK VGND VGND VPWR VPWR clknet_6_31__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26910_ _11788_ registers\[3\]\[28\] _11772_ VGND VGND VPWR VPWR _11789_ sky130_fd_sc_hd__mux2_1
X_22033_ registers\[16\]\[38\] registers\[17\]\[38\] registers\[18\]\[38\] registers\[19\]\[38\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__mux4_1
XTAP_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34019_ clknet_leaf_440_CLK _02133_ VGND VGND VPWR VPWR registers\[36\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_27890_ _12322_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26841_ net61 VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__buf_4
XTAP_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29560_ registers\[20\]\[19\] _12974_ _13222_ VGND VGND VPWR VPWR _13232_ sky130_fd_sc_hd__mux2_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26772_ registers\[40\]\[40\] _10388_ _11702_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__mux2_1
X_23984_ _10166_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28511_ _12649_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__clkbuf_1
X_25723_ registers\[48\]\[57\] _10424_ _11141_ VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29491_ _09797_ registers\[21\]\[50\] _13195_ VGND VGND VPWR VPWR _13196_ sky130_fd_sc_hd__mux2_1
X_22935_ net10 VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__clkbuf_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28442_ _11797_ registers\[28\]\[32\] _12610_ VGND VGND VPWR VPWR _12613_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25654_ registers\[48\]\[24\] _10355_ _11108_ VGND VGND VPWR VPWR _11113_ sky130_fd_sc_hd__mux2_1
X_22866_ registers\[24\]\[63\] registers\[25\]\[63\] registers\[26\]\[63\] registers\[27\]\[63\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__mux4_1
XFILLER_3_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24605_ _09535_ registers\[55\]\[10\] _10525_ VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__mux2_1
XFILLER_231_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28373_ _10014_ _10729_ VGND VGND VPWR VPWR _12576_ sky130_fd_sc_hd__nand2_8
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21817_ _08267_ _08482_ _08483_ _08270_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__a22o_1
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25585_ registers\[4\]\[57\] _10424_ _11067_ VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__mux2_1
XFILLER_71_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22797_ _07385_ _09433_ _09434_ _07395_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__a22o_1
XFILLER_197_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27324_ registers\[36\]\[15\] _10336_ _12018_ VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__mux2_1
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24536_ _09605_ registers\[56\]\[43\] _10484_ VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__mux2_1
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21748_ _08412_ _08415_ _08416_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__o21ba_1
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27255_ _11987_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24467_ _09535_ registers\[56\]\[10\] _10451_ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__mux2_1
XFILLER_200_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21679_ registers\[24\]\[28\] registers\[25\]\[28\] registers\[26\]\[28\] registers\[27\]\[28\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__mux4_1
XFILLER_123_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26206_ _10791_ registers\[44\]\[29\] _11394_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__mux2_1
XFILLER_8_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23418_ _09863_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27186_ _11951_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__clkbuf_1
X_24398_ registers\[57\]\[49\] _10407_ _10389_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26137_ _11367_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23349_ _09827_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26068_ _11331_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17910_ registers\[36\]\[52\] registers\[37\]\[52\] registers\[38\]\[52\] registers\[39\]\[52\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__mux4_1
X_25019_ net64 VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__buf_4
XFILLER_238_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1603 _14564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1614 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18890_ _05635_ _05638_ _05508_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1625 _15845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1636 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17841_ _04548_ _04616_ _04617_ _04552_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a22o_1
XANTENNA_1647 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29827_ _13372_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__clkbuf_1
XTAP_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1658 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1669 _00047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17772_ registers\[52\]\[48\] registers\[53\]\[48\] registers\[54\]\[48\] registers\[55\]\[48\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__mux4_1
X_29758_ registers\[1\]\[49\] _13037_ _13326_ VGND VGND VPWR VPWR _13336_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19511_ registers\[60\]\[32\] registers\[61\]\[32\] registers\[62\]\[32\] registers\[63\]\[32\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__mux4_1
XFILLER_43_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16723_ registers\[4\]\[18\] registers\[5\]\[18\] registers\[6\]\[18\] registers\[7\]\[18\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15219_ sky130_fd_sc_hd__mux4_1
X_28709_ _12753_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29689_ registers\[1\]\[16\] _12968_ _13293_ VGND VGND VPWR VPWR _13300_ sky130_fd_sc_hd__mux2_1
XFILLER_47_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19442_ registers\[0\]\[30\] registers\[1\]\[30\] registers\[2\]\[30\] registers\[3\]\[30\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__mux4_1
X_16654_ _14594_ VGND VGND VPWR VPWR _15152_ sky130_fd_sc_hd__buf_4
X_31720_ _14368_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_4_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31651_ _14276_ VGND VGND VPWR VPWR _14332_ sky130_fd_sc_hd__buf_6
XFILLER_222_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19373_ registers\[12\]\[28\] registers\[13\]\[28\] registers\[14\]\[28\] registers\[15\]\[28\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__mux4_1
X_16585_ registers\[16\]\[14\] registers\[17\]\[14\] registers\[18\]\[14\] registers\[19\]\[14\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _15085_ sky130_fd_sc_hd__mux4_1
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30602_ registers\[12\]\[0\] _12931_ _13780_ VGND VGND VPWR VPWR _13781_ sky130_fd_sc_hd__mux2_1
XFILLER_203_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18324_ _05077_ _05082_ _05085_ _05086_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a22o_1
XFILLER_241_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34370_ clknet_leaf_205_CLK _02484_ VGND VGND VPWR VPWR registers\[31\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31582_ registers\[63\]\[17\] net9 _14288_ VGND VGND VPWR VPWR _14296_ sky130_fd_sc_hd__mux2_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18255_ registers\[60\]\[63\] registers\[61\]\[63\] registers\[62\]\[63\] registers\[63\]\[63\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__mux4_1
X_33321_ clknet_leaf_60_CLK _01435_ VGND VGND VPWR VPWR registers\[47\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_30533_ _13744_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17206_ _15684_ _15685_ _15686_ _15687_ VGND VGND VPWR VPWR _15688_ sky130_fd_sc_hd__a22o_1
X_36040_ clknet_leaf_178_CLK _04154_ VGND VGND VPWR VPWR registers\[63\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30464_ _13707_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__clkbuf_1
X_18186_ registers\[32\]\[61\] registers\[33\]\[61\] registers\[34\]\[61\] registers\[35\]\[61\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__mux4_1
X_33252_ clknet_leaf_440_CLK _01366_ VGND VGND VPWR VPWR registers\[48\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32203_ clknet_leaf_382_CLK _00317_ VGND VGND VPWR VPWR registers\[9\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_17137_ _14555_ VGND VGND VPWR VPWR _15621_ sky130_fd_sc_hd__clkbuf_4
X_33183_ clknet_leaf_480_CLK _01297_ VGND VGND VPWR VPWR registers\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30395_ _09753_ registers\[14\]\[30\] _13671_ VGND VGND VPWR VPWR _13672_ sky130_fd_sc_hd__mux2_1
X_32134_ clknet_leaf_460_CLK _00051_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17068_ _15549_ _15551_ _15552_ _15553_ VGND VGND VPWR VPWR _15554_ sky130_fd_sc_hd__a22o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16019_ registers\[56\]\[0\] registers\[57\]\[0\] registers\[58\]\[0\] registers\[59\]\[0\]
+ _14530_ _14532_ VGND VGND VPWR VPWR _14533_ sky130_fd_sc_hd__mux4_1
XFILLER_100_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32065_ clknet_leaf_201_CLK _00243_ VGND VGND VPWR VPWR registers\[62\]\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31016_ _13998_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__clkbuf_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35824_ clknet_leaf_376_CLK _03938_ VGND VGND VPWR VPWR registers\[8\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19709_ _05080_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__buf_4
X_35755_ clknet_leaf_459_CLK _03869_ VGND VGND VPWR VPWR registers\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32967_ clknet_leaf_196_CLK _01081_ VGND VGND VPWR VPWR registers\[53\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20981_ _07671_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22720_ registers\[20\]\[58\] registers\[21\]\[58\] registers\[22\]\[58\] registers\[23\]\[58\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__mux4_1
X_34706_ clknet_leaf_96_CLK _02820_ VGND VGND VPWR VPWR registers\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31918_ _14472_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35686_ clknet_leaf_461_CLK _03800_ VGND VGND VPWR VPWR registers\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32898_ clknet_leaf_265_CLK _01012_ VGND VGND VPWR VPWR registers\[54\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34637_ clknet_leaf_148_CLK _02751_ VGND VGND VPWR VPWR registers\[27\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_22651_ _07276_ _09292_ _09293_ _07286_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__a22o_1
XFILLER_213_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31849_ _14436_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21602_ _07366_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__buf_4
XFILLER_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25370_ _10960_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__clkbuf_1
X_34568_ clknet_leaf_213_CLK _02682_ VGND VGND VPWR VPWR registers\[28\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_22582_ _07326_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__buf_6
XFILLER_146_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24321_ registers\[57\]\[24\] _10355_ _10347_ VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__mux2_1
XFILLER_166_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21533_ _07929_ _08206_ _08207_ _07932_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__a22o_1
X_33519_ clknet_leaf_361_CLK _01633_ VGND VGND VPWR VPWR registers\[44\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_34499_ clknet_leaf_225_CLK _02613_ VGND VGND VPWR VPWR registers\[2\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27040_ _11874_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_1
X_24252_ net23 VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__clkbuf_4
X_21464_ _07924_ _08139_ _08140_ _07927_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__a22o_1
XFILLER_193_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23203_ _09732_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
X_20415_ _07116_ _07119_ _06866_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__o21ba_1
X_36169_ clknet_leaf_208_CLK _04283_ VGND VGND VPWR VPWR registers\[49\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21395_ _08069_ _08072_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__o21ba_1
X_24183_ _10271_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23134_ registers\[39\]\[15\] _09689_ _09679_ VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__mux2_1
X_20346_ registers\[52\]\[56\] registers\[53\]\[56\] registers\[54\]\[56\] registers\[55\]\[56\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__mux4_1
XFILLER_88_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28991_ _12901_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__clkbuf_1
XTAP_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23065_ net57 VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__clkbuf_4
X_20277_ _06982_ _06985_ _06847_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__o21ba_1
XTAP_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27942_ registers\[32\]\[51\] _10412_ _12348_ VGND VGND VPWR VPWR _12350_ sky130_fd_sc_hd__mux2_1
XTAP_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22016_ _07324_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__clkbuf_4
XTAP_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27873_ _12313_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29612_ _13259_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__clkbuf_1
X_26824_ _11728_ registers\[3\]\[0\] _11730_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__mux2_1
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29543_ _13223_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__clkbuf_1
X_26755_ registers\[40\]\[32\] _10372_ _11691_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__mux2_1
X_23967_ _10156_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25706_ registers\[48\]\[49\] _10407_ _11130_ VGND VGND VPWR VPWR _11140_ sky130_fd_sc_hd__mux2_1
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22918_ _09540_ registers\[62\]\[12\] _09536_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__mux2_1
XFILLER_56_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26686_ _11656_ VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__buf_12
X_29474_ _09780_ registers\[21\]\[42\] _13184_ VGND VGND VPWR VPWR _13187_ sky130_fd_sc_hd__mux2_1
XFILLER_17_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23898_ _10120_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28425_ _11780_ registers\[28\]\[24\] _12599_ VGND VGND VPWR VPWR _12604_ sky130_fd_sc_hd__mux2_1
X_25637_ registers\[48\]\[16\] _10338_ _11097_ VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__mux2_1
XFILLER_232_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22849_ registers\[36\]\[63\] registers\[37\]\[63\] registers\[38\]\[63\] registers\[39\]\[63\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__mux4_1
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28356_ _12567_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__clkbuf_1
X_16370_ registers\[4\]\[8\] registers\[5\]\[8\] registers\[6\]\[8\] registers\[7\]\[8\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _14876_ sky130_fd_sc_hd__mux4_1
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25568_ registers\[4\]\[49\] _10407_ _11056_ VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__mux2_1
XFILLER_13_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27307_ registers\[36\]\[7\] _10319_ _12007_ VGND VGND VPWR VPWR _12015_ sky130_fd_sc_hd__mux2_1
XFILLER_158_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24519_ _09588_ registers\[56\]\[35\] _10473_ VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__mux2_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28287_ _12531_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__clkbuf_1
X_25499_ registers\[4\]\[16\] _10338_ _11023_ VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__mux2_1
XFILLER_200_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18040_ _04683_ _04809_ _04810_ _04686_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__a22o_1
X_27238_ _11978_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27169_ _11942_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30180_ registers\[16\]\[57\] _13054_ _13550_ VGND VGND VPWR VPWR _13558_ sky130_fd_sc_hd__mux2_1
XFILLER_99_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19991_ registers\[56\]\[46\] registers\[57\]\[46\] registers\[58\]\[46\] registers\[59\]\[46\]
+ _06644_ _06434_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux4_1
XFILLER_180_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18942_ registers\[8\]\[16\] registers\[9\]\[16\] registers\[10\]\[16\] registers\[11\]\[16\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__mux4_1
XANTENNA_1400 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1411 _00179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1422 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1433 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18873_ _05412_ _05620_ _05621_ _05416_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__a22o_1
XFILLER_239_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1444 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1455 _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1466 _05162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17824_ _04580_ _04587_ _04594_ _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__or4_2
XANTENNA_1477 _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33870_ clknet_leaf_134_CLK _01984_ VGND VGND VPWR VPWR registers\[38\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1488 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1499 _07328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32821_ clknet_leaf_353_CLK _00935_ VGND VGND VPWR VPWR registers\[55\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_17755_ registers\[32\]\[48\] registers\[33\]\[48\] registers\[34\]\[48\] registers\[35\]\[48\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__mux4_1
X_35540_ clknet_leaf_81_CLK _03654_ VGND VGND VPWR VPWR registers\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_16706_ _14496_ VGND VGND VPWR VPWR _15202_ sky130_fd_sc_hd__clkbuf_4
X_32752_ clknet_leaf_366_CLK _00866_ VGND VGND VPWR VPWR registers\[56\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17686_ _04333_ _04465_ _04466_ _04338_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a22o_1
XFILLER_208_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31703_ registers\[59\]\[10\] net2 _14359_ VGND VGND VPWR VPWR _14360_ sky130_fd_sc_hd__mux2_1
X_19425_ registers\[44\]\[30\] registers\[45\]\[30\] registers\[46\]\[30\] registers\[47\]\[30\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux4_2
X_35471_ clknet_leaf_140_CLK _03585_ VGND VGND VPWR VPWR registers\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16637_ _14548_ VGND VGND VPWR VPWR _15135_ sky130_fd_sc_hd__buf_4
X_32683_ clknet_leaf_424_CLK _00797_ VGND VGND VPWR VPWR registers\[57\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34422_ clknet_leaf_426_CLK _02536_ VGND VGND VPWR VPWR registers\[30\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_19356_ _05080_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__buf_6
X_31634_ _14323_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16568_ registers\[48\]\[14\] registers\[49\]\[14\] registers\[50\]\[14\] registers\[51\]\[14\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15068_ sky130_fd_sc_hd__mux4_1
XFILLER_210_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18307_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__buf_4
XFILLER_52_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34353_ clknet_leaf_386_CLK _02467_ VGND VGND VPWR VPWR registers\[31\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31565_ registers\[63\]\[9\] net64 _14277_ VGND VGND VPWR VPWR _14287_ sky130_fd_sc_hd__mux2_1
X_19287_ _05747_ _06022_ _06023_ _05753_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__a22o_1
X_16499_ _14581_ VGND VGND VPWR VPWR _15001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33304_ clknet_leaf_31_CLK _01418_ VGND VGND VPWR VPWR registers\[47\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_18238_ _14558_ _05001_ _05002_ _14568_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__a22o_1
X_30516_ _13735_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34284_ clknet_leaf_325_CLK _02398_ VGND VGND VPWR VPWR registers\[32\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_31496_ _09775_ registers\[6\]\[40\] _14250_ VGND VGND VPWR VPWR _14251_ sky130_fd_sc_hd__mux2_1
XFILLER_209_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36023_ clknet_leaf_330_CLK _04137_ VGND VGND VPWR VPWR registers\[63\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_30447_ _09808_ registers\[14\]\[55\] _13693_ VGND VGND VPWR VPWR _13699_ sky130_fd_sc_hd__mux2_1
X_33235_ clknet_leaf_70_CLK _01349_ VGND VGND VPWR VPWR registers\[48\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18169_ registers\[8\]\[60\] registers\[9\]\[60\] registers\[10\]\[60\] registers\[11\]\[60\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux4_1
XFILLER_198_1079 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20200_ _06911_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21180_ _07586_ _07863_ _07864_ _07589_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__a22o_1
X_33166_ clknet_leaf_139_CLK _01280_ VGND VGND VPWR VPWR registers\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_30378_ _09717_ registers\[14\]\[22\] _13660_ VGND VGND VPWR VPWR _13663_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20131_ registers\[44\]\[50\] registers\[45\]\[50\] registers\[46\]\[50\] registers\[47\]\[50\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux4_1
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32117_ clknet_leaf_467_CLK _00032_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dfxtp_1
X_33097_ clknet_leaf_207_CLK _01211_ VGND VGND VPWR VPWR registers\[51\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20062_ _05080_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__clkbuf_4
X_32048_ clknet_leaf_371_CLK _00226_ VGND VGND VPWR VPWR registers\[62\]\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24870_ _09529_ registers\[53\]\[7\] _10658_ VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__mux2_1
XFILLER_112_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23821_ _10079_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__clkbuf_1
X_35807_ clknet_leaf_484_CLK _03921_ VGND VGND VPWR VPWR registers\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33999_ clknet_leaf_133_CLK _02113_ VGND VGND VPWR VPWR registers\[36\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26540_ _11579_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23752_ _10043_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
X_35738_ clknet_leaf_479_CLK _03852_ VGND VGND VPWR VPWR registers\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_308 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20964_ registers\[8\]\[8\] registers\[9\]\[8\] registers\[10\]\[8\] registers\[11\]\[8\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__mux4_1
XANTENNA_319 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ registers\[48\]\[58\] registers\[49\]\[58\] registers\[50\]\[58\] registers\[51\]\[58\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__mux4_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26471_ _11543_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__clkbuf_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23683_ _10005_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
X_35669_ clknet_leaf_79_CLK _03783_ VGND VGND VPWR VPWR registers\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ registers\[4\]\[6\] registers\[5\]\[6\] registers\[6\]\[6\] registers\[7\]\[6\]
+ _07362_ _07364_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28210_ _11834_ registers\[30\]\[50\] _12490_ VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__mux2_1
XFILLER_148_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25422_ _10987_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22634_ _09277_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
X_29190_ _13028_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_224_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28141_ _12454_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25353_ _10951_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22565_ registers\[28\]\[53\] registers\[29\]\[53\] registers\[30\]\[53\] registers\[31\]\[53\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24304_ net11 VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__buf_4
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28072_ _11832_ registers\[31\]\[49\] _12408_ VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21516_ registers\[36\]\[24\] registers\[37\]\[24\] registers\[38\]\[24\] registers\[39\]\[24\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25284_ _10914_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__clkbuf_1
X_22496_ registers\[20\]\[51\] registers\[21\]\[51\] registers\[22\]\[51\] registers\[23\]\[51\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__mux4_1
XFILLER_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27023_ _11728_ registers\[38\]\[0\] _11865_ VGND VGND VPWR VPWR _11866_ sky130_fd_sc_hd__mux2_1
XFILLER_181_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24235_ _10298_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21447_ _07285_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24166_ _10262_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21378_ registers\[48\]\[20\] registers\[49\]\[20\] registers\[50\]\[20\] registers\[51\]\[20\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__mux4_1
X_23117_ net2 VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__clkbuf_8
XFILLER_79_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20329_ registers\[28\]\[55\] registers\[29\]\[55\] registers\[30\]\[55\] registers\[31\]\[55\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__mux4_1
X_24097_ _10225_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
X_28974_ _12892_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23048_ _09628_ registers\[62\]\[54\] _09620_ VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__mux2_1
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27925_ registers\[32\]\[43\] _10395_ _12337_ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__mux2_1
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27856_ registers\[32\]\[10\] _10325_ _12304_ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__mux2_1
XFILLER_237_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26807_ registers\[40\]\[57\] _10424_ _11713_ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__mux2_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24999_ _10735_ registers\[52\]\[2\] _10731_ VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__mux2_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27787_ _12268_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__clkbuf_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29526_ _13214_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__clkbuf_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ registers\[16\]\[41\] registers\[17\]\[41\] registers\[18\]\[41\] registers\[19\]\[41\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__mux4_1
XFILLER_57_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26738_ registers\[40\]\[24\] _10355_ _11680_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__mux2_1
XFILLER_217_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_820 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_831 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_842 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17471_ _15924_ _15931_ _15938_ _15945_ VGND VGND VPWR VPWR _15946_ sky130_fd_sc_hd__or4_1
X_26669_ _10848_ registers\[41\]\[56\] _11641_ VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__mux2_1
XFILLER_232_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29457_ _09762_ registers\[21\]\[34\] _13173_ VGND VGND VPWR VPWR _13178_ sky130_fd_sc_hd__mux2_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_853 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_864 _09335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_875 _09527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19210_ _05926_ _05933_ _05942_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__or4_4
XFILLER_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_233_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16422_ _14524_ VGND VGND VPWR VPWR _14926_ sky130_fd_sc_hd__clkbuf_4
X_28408_ _11763_ registers\[28\]\[16\] _12588_ VGND VGND VPWR VPWR _12595_ sky130_fd_sc_hd__mux2_1
XANTENNA_886 _09588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29388_ _09660_ registers\[21\]\[1\] _13140_ VGND VGND VPWR VPWR _13142_ sky130_fd_sc_hd__mux2_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_897 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16353_ _14496_ VGND VGND VPWR VPWR _14859_ sky130_fd_sc_hd__clkbuf_4
X_19141_ _05882_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28339_ _12558_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19072_ registers\[44\]\[20\] registers\[45\]\[20\] registers\[46\]\[20\] registers\[47\]\[20\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__mux4_2
X_31350_ registers\[7\]\[35\] net29 _14168_ VGND VGND VPWR VPWR _14174_ sky130_fd_sc_hd__mux2_1
XFILLER_173_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16284_ _14548_ VGND VGND VPWR VPWR _14792_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_970 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30301_ registers\[15\]\[50\] _13039_ _13621_ VGND VGND VPWR VPWR _13622_ sky130_fd_sc_hd__mux2_1
X_18023_ registers\[4\]\[55\] registers\[5\]\[55\] registers\[6\]\[55\] registers\[7\]\[55\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__mux4_1
X_31281_ registers\[7\]\[2\] net23 _14135_ VGND VGND VPWR VPWR _14138_ sky130_fd_sc_hd__mux2_1
XFILLER_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_246_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33020_ clknet_leaf_290_CLK _01134_ VGND VGND VPWR VPWR registers\[52\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_30232_ _13585_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30163_ registers\[16\]\[49\] _13037_ _13539_ VGND VGND VPWR VPWR _13549_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19974_ _06688_ _06691_ _06523_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18925_ registers\[40\]\[16\] registers\[41\]\[16\] registers\[42\]\[16\] registers\[43\]\[16\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__mux4_1
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34971_ clknet_leaf_490_CLK _03085_ VGND VGND VPWR VPWR registers\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_30094_ registers\[16\]\[16\] _12968_ _13506_ VGND VGND VPWR VPWR _13513_ sky130_fd_sc_hd__mux2_1
XANTENNA_1230 _00034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1241 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1252 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_295_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_295_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33922_ clknet_leaf_261_CLK _02036_ VGND VGND VPWR VPWR registers\[38\]\[52\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1263 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18856_ _05602_ _05605_ _05508_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__o21ba_1
XTAP_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1274 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1285 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1296 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17807_ registers\[52\]\[49\] registers\[53\]\[49\] registers\[54\]\[49\] registers\[55\]\[49\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__mux4_1
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33853_ clknet_leaf_299_CLK _01967_ VGND VGND VPWR VPWR registers\[3\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18787_ _05517_ _05524_ _05531_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__or4_2
X_15999_ _14504_ VGND VGND VPWR VPWR _14513_ sky130_fd_sc_hd__clkbuf_4
XFILLER_212_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32804_ clknet_leaf_442_CLK _00918_ VGND VGND VPWR VPWR registers\[55\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_17738_ registers\[8\]\[47\] registers\[9\]\[47\] registers\[10\]\[47\] registers\[11\]\[47\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__mux4_1
XFILLER_209_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33784_ clknet_leaf_340_CLK _01898_ VGND VGND VPWR VPWR registers\[40\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_30996_ _13987_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35523_ clknet_leaf_239_CLK _03637_ VGND VGND VPWR VPWR registers\[13\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_32735_ clknet_leaf_38_CLK _00849_ VGND VGND VPWR VPWR registers\[56\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17669_ registers\[0\]\[45\] registers\[1\]\[45\] registers\[2\]\[45\] registers\[3\]\[45\]
+ _15967_ _15968_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_1209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19408_ registers\[4\]\[29\] registers\[5\]\[29\] registers\[6\]\[29\] registers\[7\]\[29\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__mux4_1
XFILLER_39_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35454_ clknet_leaf_196_CLK _03568_ VGND VGND VPWR VPWR registers\[14\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20680_ _07316_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__buf_12
X_32666_ clknet_leaf_84_CLK _00780_ VGND VGND VPWR VPWR registers\[57\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34405_ clknet_leaf_464_CLK _02519_ VGND VGND VPWR VPWR registers\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31617_ _14314_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__clkbuf_1
X_19339_ registers\[24\]\[27\] registers\[25\]\[27\] registers\[26\]\[27\] registers\[27\]\[27\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__mux4_1
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35385_ clknet_leaf_303_CLK _03499_ VGND VGND VPWR VPWR registers\[15\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_32597_ clknet_leaf_71_CLK _00711_ VGND VGND VPWR VPWR registers\[58\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22350_ _08766_ _09000_ _09001_ _08771_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__a22o_1
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34336_ clknet_leaf_488_CLK _02450_ VGND VGND VPWR VPWR registers\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31548_ _14278_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21301_ _07978_ _07981_ _07711_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__o21ba_1
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22281_ _08931_ _08934_ _08773_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__o21ba_1
X_34267_ clknet_leaf_18_CLK _02381_ VGND VGND VPWR VPWR registers\[32\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31479_ _09758_ registers\[6\]\[32\] _14239_ VGND VGND VPWR VPWR _14242_ sky130_fd_sc_hd__mux2_1
XFILLER_117_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24020_ _10185_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
X_36006_ clknet_leaf_450_CLK _04120_ VGND VGND VPWR VPWR registers\[63\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33218_ clknet_leaf_234_CLK _01332_ VGND VGND VPWR VPWR registers\[4\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_21232_ registers\[56\]\[16\] registers\[57\]\[16\] registers\[58\]\[16\] registers\[59\]\[16\]
+ _07851_ _07641_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__mux4_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34198_ clknet_leaf_122_CLK _02312_ VGND VGND VPWR VPWR registers\[33\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33149_ clknet_leaf_290_CLK _01263_ VGND VGND VPWR VPWR registers\[50\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_21163_ registers\[36\]\[14\] registers\[37\]\[14\] registers\[38\]\[14\] registers\[39\]\[14\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__mux4_1
XFILLER_160_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20114_ registers\[4\]\[49\] registers\[5\]\[49\] registers\[6\]\[49\] registers\[7\]\[49\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux4_1
X_25971_ _11280_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
X_21094_ _07352_ VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_286_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_286_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27710_ registers\[33\]\[5\] _10315_ _12222_ VGND VGND VPWR VPWR _12228_ sky130_fd_sc_hd__mux2_1
X_20045_ registers\[24\]\[47\] registers\[25\]\[47\] registers\[26\]\[47\] registers\[27\]\[47\]
+ _06660_ _06661_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__mux4_1
XFILLER_24_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24922_ _10693_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28690_ _12743_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24853_ _10656_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27641_ _12191_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_949 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23804_ _10070_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27572_ _12155_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__clkbuf_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24784_ _09577_ registers\[54\]\[30\] _10620_ VGND VGND VPWR VPWR _10621_ sky130_fd_sc_hd__mux2_1
XANTENNA_105 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21996_ registers\[20\]\[37\] registers\[21\]\[37\] registers\[22\]\[37\] registers\[23\]\[37\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__mux4_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26523_ _10838_ registers\[42\]\[51\] _11569_ VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__mux2_1
XANTENNA_127 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29311_ _09751_ registers\[22\]\[29\] _13091_ VGND VGND VPWR VPWR _13101_ sky130_fd_sc_hd__mux2_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23735_ _10034_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _07440_ _07636_ _07637_ _07443_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__a22o_1
XANTENNA_149 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29242_ _13063_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26454_ _11534_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_1
X_23666_ _09996_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__clkbuf_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _07567_ _07570_ _07310_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__o21ba_1
XFILLER_214_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25405_ _10978_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__clkbuf_1
X_22617_ _09020_ _09259_ _09260_ _09024_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__a22o_1
X_29173_ registers\[23\]\[39\] _13016_ _12998_ VGND VGND VPWR VPWR _13017_ sky130_fd_sc_hd__mux2_1
X_26385_ _11442_ VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__buf_6
XFILLER_139_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23597_ _09960_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_210_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_210_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28124_ _12445_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__clkbuf_1
X_25336_ _10942_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__clkbuf_1
X_22548_ _09012_ _09192_ _09193_ _09018_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__a22o_1
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_9_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_9_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_182_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28055_ _12409_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__clkbuf_1
X_25267_ _10905_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__clkbuf_1
X_22479_ registers\[48\]\[51\] registers\[49\]\[51\] registers\[50\]\[51\] registers\[51\]\[51\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__mux4_1
X_27006_ _11853_ registers\[3\]\[59\] _11835_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__mux2_1
X_24218_ _09622_ registers\[58\]\[51\] _10288_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__mux2_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25198_ _10869_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24149_ _10253_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16971_ _15290_ _15458_ _15459_ _15293_ VGND VGND VPWR VPWR _15460_ sky130_fd_sc_hd__a22o_1
X_28957_ registers\[24\]\[20\] _10346_ _12883_ VGND VGND VPWR VPWR _12884_ sky130_fd_sc_hd__mux2_1
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_277_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_277_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18710_ _05150_ _05462_ _05463_ _05160_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__a22o_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27908_ registers\[32\]\[35\] _10378_ _12326_ VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__mux2_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _06379_ _06414_ _06415_ _06382_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a22o_1
X_28888_ _12847_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__clkbuf_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _05396_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27839_ registers\[32\]\[2\] _10309_ _12293_ VGND VGND VPWR VPWR _12296_ sky130_fd_sc_hd__mux2_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30850_ _09806_ registers\[11\]\[54\] _13906_ VGND VGND VPWR VPWR _13911_ sky130_fd_sc_hd__mux2_1
X_18572_ registers\[40\]\[6\] registers\[41\]\[6\] registers\[42\]\[6\] registers\[43\]\[6\]
+ _05198_ _05199_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__mux4_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29509_ _09817_ registers\[21\]\[59\] _13195_ VGND VGND VPWR VPWR _13205_ sky130_fd_sc_hd__mux2_1
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _15684_ _04307_ _04308_ _15687_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a22o_1
XFILLER_45_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30781_ _09702_ registers\[11\]\[21\] _13873_ VGND VGND VPWR VPWR _13875_ sky130_fd_sc_hd__mux2_1
XANTENNA_650 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_661 _05297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32520_ clknet_leaf_178_CLK _00634_ VGND VGND VPWR VPWR registers\[60\]\[58\] sky130_fd_sc_hd__dfxtp_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_672 _05623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17454_ registers\[52\]\[39\] registers\[53\]\[39\] registers\[54\]\[39\] registers\[55\]\[39\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _15929_ sky130_fd_sc_hd__mux4_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_683 _06171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_694 _07135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16405_ registers\[24\]\[9\] registers\[25\]\[9\] registers\[26\]\[9\] registers\[27\]\[9\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14910_ sky130_fd_sc_hd__mux4_1
X_32451_ clknet_leaf_204_CLK _00565_ VGND VGND VPWR VPWR registers\[29\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17385_ registers\[8\]\[37\] registers\[9\]\[37\] registers\[10\]\[37\] registers\[11\]\[37\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15862_ sky130_fd_sc_hd__mux4_1
XFILLER_242_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_201_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_201_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_31402_ registers\[7\]\[60\] net57 _14134_ VGND VGND VPWR VPWR _14201_ sky130_fd_sc_hd__mux2_1
XFILLER_13_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19124_ _05755_ _05864_ _05865_ _05759_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a22o_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16336_ registers\[28\]\[7\] registers\[29\]\[7\] registers\[30\]\[7\] registers\[31\]\[7\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14843_ sky130_fd_sc_hd__mux4_1
XFILLER_125_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35170_ clknet_leaf_474_CLK _03284_ VGND VGND VPWR VPWR registers\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_32382_ clknet_leaf_293_CLK _00496_ VGND VGND VPWR VPWR registers\[61\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34121_ clknet_leaf_237_CLK _02235_ VGND VGND VPWR VPWR registers\[35\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16267_ registers\[20\]\[5\] registers\[21\]\[5\] registers\[22\]\[5\] registers\[23\]\[5\]
+ _14606_ _14608_ VGND VGND VPWR VPWR _14776_ sky130_fd_sc_hd__mux4_1
X_19055_ registers\[4\]\[19\] registers\[5\]\[19\] registers\[6\]\[19\] registers\[7\]\[19\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__mux4_1
X_31333_ registers\[7\]\[27\] net20 _14157_ VGND VGND VPWR VPWR _14165_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18006_ registers\[32\]\[55\] registers\[33\]\[55\] registers\[34\]\[55\] registers\[35\]\[55\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__mux4_1
XFILLER_127_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34052_ clknet_leaf_252_CLK _02166_ VGND VGND VPWR VPWR registers\[36\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31264_ _14128_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__clkbuf_1
X_16198_ registers\[16\]\[3\] registers\[17\]\[3\] registers\[18\]\[3\] registers\[19\]\[3\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14709_ sky130_fd_sc_hd__mux4_1
XFILLER_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33003_ clknet_leaf_420_CLK _01117_ VGND VGND VPWR VPWR registers\[52\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_30215_ _13576_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31195_ _14092_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30146_ _13540_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19957_ _06576_ _06673_ _06674_ _06579_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__a22o_1
XFILLER_141_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_268_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_268_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18908_ _05053_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__clkbuf_4
X_34954_ clknet_leaf_143_CLK _03068_ VGND VGND VPWR VPWR registers\[22\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_30077_ registers\[16\]\[8\] _12951_ _13495_ VGND VGND VPWR VPWR _13504_ sky130_fd_sc_hd__mux2_1
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19888_ _06569_ _06606_ _06607_ _06574_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__a22o_1
XANTENNA_1060 _13850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1071 _14347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33905_ clknet_leaf_359_CLK _02019_ VGND VGND VPWR VPWR registers\[38\]\[35\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1082 _14496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1093 _14524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18839_ _05412_ _05587_ _05588_ _05416_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a22o_1
XFILLER_28_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34885_ clknet_leaf_212_CLK _02999_ VGND VGND VPWR VPWR registers\[23\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33836_ clknet_leaf_388_CLK _01950_ VGND VGND VPWR VPWR registers\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_21850_ _07303_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__buf_6
XFILLER_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20801_ registers\[20\]\[3\] registers\[21\]\[3\] registers\[22\]\[3\] registers\[23\]\[3\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__mux4_1
XFILLER_184_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21781_ _08267_ _08447_ _08448_ _08270_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__a22o_1
XFILLER_35_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33767_ clknet_leaf_430_CLK _01881_ VGND VGND VPWR VPWR registers\[40\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_30979_ registers\[10\]\[51\] _13042_ _13977_ VGND VGND VPWR VPWR _13979_ sky130_fd_sc_hd__mux2_1
XFILLER_212_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23520_ _09607_ registers\[19\]\[44\] _09914_ VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__mux2_1
X_35506_ clknet_leaf_356_CLK _03620_ VGND VGND VPWR VPWR registers\[13\]\[36\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_440_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_440_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20732_ _07386_ _07428_ _07429_ _07396_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__a22o_1
X_32718_ clknet_leaf_173_CLK _00832_ VGND VGND VPWR VPWR registers\[56\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33698_ clknet_leaf_56_CLK _01812_ VGND VGND VPWR VPWR registers\[41\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35437_ clknet_leaf_393_CLK _03551_ VGND VGND VPWR VPWR registers\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23451_ _09538_ registers\[19\]\[11\] _09881_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__mux2_1
X_20663_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__buf_6
X_32649_ clknet_leaf_209_CLK _00763_ VGND VGND VPWR VPWR registers\[58\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_22402_ _09048_ _09051_ _08740_ VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__o21ba_1
XFILLER_195_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26170_ _11385_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
X_23382_ registers\[39\]\[44\] _09784_ _09840_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__mux2_1
X_35368_ clknet_leaf_399_CLK _03482_ VGND VGND VPWR VPWR registers\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20594_ net73 net74 VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__and2_1
XFILLER_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25121_ _10818_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__clkbuf_1
X_34319_ clknet_leaf_110_CLK _02433_ VGND VGND VPWR VPWR registers\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_22333_ _08669_ _08983_ _08984_ _08675_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__a22o_1
XFILLER_191_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35299_ clknet_leaf_474_CLK _03413_ VGND VGND VPWR VPWR registers\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25052_ _10771_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
X_22264_ _08677_ _08916_ _08917_ _08681_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__a22o_1
XFILLER_105_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24003_ _10176_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21215_ _07895_ _07898_ _07730_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__o21ba_2
X_29860_ registers\[18\]\[33\] _13004_ _13386_ VGND VGND VPWR VPWR _13390_ sky130_fd_sc_hd__mux2_1
X_22195_ _08669_ _08849_ _08850_ _08675_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__a22o_1
XFILLER_160_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28811_ _11761_ registers\[25\]\[15\] _12801_ VGND VGND VPWR VPWR _12807_ sky130_fd_sc_hd__mux2_1
X_21146_ registers\[12\]\[13\] registers\[13\]\[13\] registers\[14\]\[13\] registers\[15\]\[13\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__mux4_1
X_29791_ registers\[18\]\[0\] _12931_ _13353_ VGND VGND VPWR VPWR _13354_ sky130_fd_sc_hd__mux2_1
XFILLER_63_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_259_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_259_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_1333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28742_ _12770_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__clkbuf_1
X_21077_ registers\[4\]\[11\] registers\[5\]\[11\] registers\[6\]\[11\] registers\[7\]\[11\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__mux4_1
X_25954_ _11271_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20028_ registers\[36\]\[47\] registers\[37\]\[47\] registers\[38\]\[47\] registers\[39\]\[47\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__mux4_1
X_24905_ _10684_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
X_25885_ _11235_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
X_28673_ _12734_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27624_ _12182_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__clkbuf_1
X_24836_ _09630_ registers\[54\]\[55\] _10642_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__mux2_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27555_ _11857_ registers\[35\]\[61\] _12077_ VGND VGND VPWR VPWR _12145_ sky130_fd_sc_hd__mux2_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24767_ _09561_ registers\[54\]\[22\] _10609_ VGND VGND VPWR VPWR _10612_ sky130_fd_sc_hd__mux2_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ registers\[48\]\[37\] registers\[49\]\[37\] registers\[50\]\[37\] registers\[51\]\[37\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__mux4_1
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_431_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_431_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_215_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23718_ _10025_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
X_26506_ _10821_ registers\[42\]\[43\] _11558_ VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__mux2_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27486_ _11788_ registers\[35\]\[28\] _12100_ VGND VGND VPWR VPWR _12109_ sky130_fd_sc_hd__mux2_1
XFILLER_214_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24698_ _10574_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29225_ net52 VGND VGND VPWR VPWR _13052_ sky130_fd_sc_hd__clkbuf_4
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26437_ _10751_ registers\[42\]\[10\] _11525_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__mux2_1
X_23649_ registers\[61\]\[40\] _09775_ _09987_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__mux2_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17170_ _15341_ _15651_ _15652_ _15344_ VGND VGND VPWR VPWR _15653_ sky130_fd_sc_hd__a22o_1
X_29156_ _13005_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__clkbuf_1
X_26368_ _11489_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16121_ registers\[0\]\[1\] registers\[1\]\[1\] registers\[2\]\[1\] registers\[3\]\[1\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14634_ sky130_fd_sc_hd__mux4_1
X_28107_ _11732_ registers\[30\]\[1\] _12435_ VGND VGND VPWR VPWR _12437_ sky130_fd_sc_hd__mux2_1
X_25319_ _10932_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26299_ _10749_ registers\[43\]\[9\] _11443_ VGND VGND VPWR VPWR _11453_ sky130_fd_sc_hd__mux2_1
XFILLER_127_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29087_ registers\[23\]\[11\] _12958_ _12956_ VGND VGND VPWR VPWR _12959_ sky130_fd_sc_hd__mux2_1
XFILLER_194_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16052_ registers\[0\]\[0\] registers\[1\]\[0\] registers\[2\]\[0\] registers\[3\]\[0\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14566_ sky130_fd_sc_hd__mux4_1
X_28038_ _12400_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30000_ _13463_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19811_ registers\[20\]\[40\] registers\[21\]\[40\] registers\[22\]\[40\] registers\[23\]\[40\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__mux4_1
XFILLER_29_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29989_ registers\[17\]\[30\] _12997_ _13457_ VGND VGND VPWR VPWR _13458_ sky130_fd_sc_hd__mux2_1
XFILLER_96_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19742_ _05067_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__buf_4
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16954_ registers\[48\]\[25\] registers\[49\]\[25\] registers\[50\]\[25\] registers\[51\]\[25\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15443_ sky130_fd_sc_hd__mux4_1
XFILLER_96_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31951_ clknet_leaf_492_CLK _00139_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_1
X_19673_ _05120_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__buf_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16885_ _15341_ _15374_ _15375_ _15344_ VGND VGND VPWR VPWR _15376_ sky130_fd_sc_hd__a22o_1
X_18624_ _05089_ _05378_ _05379_ _05100_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__a22o_1
X_30902_ _13938_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__clkbuf_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34670_ clknet_leaf_410_CLK _02784_ VGND VGND VPWR VPWR registers\[26\]\[32\] sky130_fd_sc_hd__dfxtp_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31882_ _09756_ registers\[49\]\[31\] _14452_ VGND VGND VPWR VPWR _14454_ sky130_fd_sc_hd__mux2_1
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33621_ clknet_leaf_124_CLK _01735_ VGND VGND VPWR VPWR registers\[42\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_30833_ _09788_ registers\[11\]\[46\] _13895_ VGND VGND VPWR VPWR _13902_ sky130_fd_sc_hd__mux2_1
X_18555_ _05053_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__buf_4
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_422_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_422_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17506_ _04289_ _04290_ _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a22o_1
XFILLER_244_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33552_ clknet_leaf_129_CLK _01666_ VGND VGND VPWR VPWR registers\[43\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18486_ _05089_ _05244_ _05245_ _05100_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__a22o_1
X_30764_ _09685_ registers\[11\]\[13\] _13862_ VGND VGND VPWR VPWR _13866_ sky130_fd_sc_hd__mux2_1
XFILLER_221_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_480 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_491 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32503_ clknet_leaf_331_CLK _00617_ VGND VGND VPWR VPWR registers\[60\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17437_ _15638_ _15911_ _15912_ _15643_ VGND VGND VPWR VPWR _15913_ sky130_fd_sc_hd__a22o_1
X_33483_ clknet_leaf_165_CLK _01597_ VGND VGND VPWR VPWR registers\[45\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30695_ _13829_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_16 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35222_ clknet_leaf_89_CLK _03336_ VGND VGND VPWR VPWR registers\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_27 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32434_ clknet_leaf_412_CLK _00548_ VGND VGND VPWR VPWR registers\[29\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_49 _00046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17368_ _15845_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19107_ _05844_ _05845_ _05848_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__a22o_1
X_35153_ clknet_leaf_101_CLK _03267_ VGND VGND VPWR VPWR registers\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16319_ registers\[56\]\[7\] registers\[57\]\[7\] registers\[58\]\[7\] registers\[59\]\[7\]
+ _14723_ _14532_ VGND VGND VPWR VPWR _14826_ sky130_fd_sc_hd__mux4_1
XFILLER_174_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32365_ clknet_leaf_374_CLK _00479_ VGND VGND VPWR VPWR registers\[61\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_17299_ registers\[40\]\[35\] registers\[41\]\[35\] registers\[42\]\[35\] registers\[43\]\[35\]
+ _15678_ _15679_ VGND VGND VPWR VPWR _15778_ sky130_fd_sc_hd__mux4_1
XFILLER_88_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34104_ clknet_leaf_337_CLK _02218_ VGND VGND VPWR VPWR registers\[35\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31316_ registers\[7\]\[19\] net11 _14146_ VGND VGND VPWR VPWR _14156_ sky130_fd_sc_hd__mux2_1
X_19038_ registers\[32\]\[19\] registers\[33\]\[19\] registers\[34\]\[19\] registers\[35\]\[19\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__mux4_1
X_35084_ clknet_leaf_143_CLK _03198_ VGND VGND VPWR VPWR registers\[20\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput101 net101 VGND VGND VPWR VPWR D1[1] sky130_fd_sc_hd__buf_2
X_32296_ clknet_leaf_406_CLK _00410_ VGND VGND VPWR VPWR registers\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput112 net112 VGND VGND VPWR VPWR D1[2] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_489_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_489_CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput123 net123 VGND VGND VPWR VPWR D1[3] sky130_fd_sc_hd__buf_2
X_34035_ clknet_leaf_348_CLK _02149_ VGND VGND VPWR VPWR registers\[36\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31247_ registers\[8\]\[50\] net46 _14119_ VGND VGND VPWR VPWR _14120_ sky130_fd_sc_hd__mux2_1
Xoutput134 net134 VGND VGND VPWR VPWR D1[4] sky130_fd_sc_hd__buf_2
XFILLER_99_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput145 net145 VGND VGND VPWR VPWR D1[5] sky130_fd_sc_hd__buf_2
Xoutput156 net156 VGND VGND VPWR VPWR D2[11] sky130_fd_sc_hd__buf_2
XFILLER_86_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21000_ _07581_ _07688_ _07689_ _07584_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a22o_1
XFILLER_130_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput167 net167 VGND VGND VPWR VPWR D2[21] sky130_fd_sc_hd__buf_2
XFILLER_142_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput178 net178 VGND VGND VPWR VPWR D2[31] sky130_fd_sc_hd__buf_2
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput189 net189 VGND VGND VPWR VPWR D2[41] sky130_fd_sc_hd__buf_2
XFILLER_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31178_ _14083_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30129_ _13531_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35986_ clknet_leaf_181_CLK _04100_ VGND VGND VPWR VPWR registers\[63\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34937_ clknet_leaf_308_CLK _03051_ VGND VGND VPWR VPWR registers\[22\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_22951_ net16 VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__buf_2
XFILLER_25_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21902_ registers\[44\]\[35\] registers\[45\]\[35\] registers\[46\]\[35\] registers\[47\]\[35\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__mux4_1
X_25670_ _11121_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22882_ _09516_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
X_34868_ clknet_leaf_384_CLK _02982_ VGND VGND VPWR VPWR registers\[23\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24621_ _09552_ registers\[55\]\[18\] _10525_ VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__mux2_1
X_33819_ clknet_leaf_478_CLK _01933_ VGND VGND VPWR VPWR registers\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21833_ registers\[40\]\[33\] registers\[41\]\[33\] registers\[42\]\[33\] registers\[43\]\[33\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__mux4_1
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34799_ clknet_leaf_382_CLK _02913_ VGND VGND VPWR VPWR registers\[24\]\[33\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_413_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_413_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27340_ _12032_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__clkbuf_1
X_24552_ _10496_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21764_ _08432_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23503_ _09590_ registers\[19\]\[36\] _09903_ VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__mux2_1
XFILLER_58_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27271_ _11843_ registers\[37\]\[54\] _11991_ VGND VGND VPWR VPWR _11996_ sky130_fd_sc_hd__mux2_1
Xclkbuf_6_54__f_CLK clknet_5_27_0_CLK VGND VGND VPWR VPWR clknet_6_54__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20715_ _07313_ _07411_ _07412_ _07322_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__a22o_1
XFILLER_211_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24483_ _09552_ registers\[56\]\[18\] _10451_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__mux2_1
X_21695_ _08126_ _08363_ _08364_ _08129_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__a22o_1
XFILLER_145_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29010_ _12911_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__clkbuf_1
X_26222_ _11412_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
X_23434_ _09521_ registers\[19\]\[3\] _09870_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__mux2_1
X_20646_ _07289_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__buf_6
XFILLER_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26153_ _11376_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23365_ registers\[39\]\[36\] _09766_ _09829_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__mux2_1
X_20577_ _07275_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25104_ _10806_ registers\[52\]\[36\] _10794_ VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__mux2_1
X_22316_ registers\[28\]\[46\] registers\[29\]\[46\] registers\[30\]\[46\] registers\[31\]\[46\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__mux4_1
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26084_ _10804_ registers\[45\]\[35\] _11334_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__mux2_1
X_23296_ _09792_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
X_29912_ registers\[18\]\[58\] _13056_ _13408_ VGND VGND VPWR VPWR _13417_ sky130_fd_sc_hd__mux2_1
X_25035_ net6 VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__clkbuf_4
X_22247_ registers\[20\]\[44\] registers\[21\]\[44\] registers\[22\]\[44\] registers\[23\]\[44\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__mux4_1
XFILLER_156_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_913 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29843_ registers\[18\]\[25\] _12987_ _13375_ VGND VGND VPWR VPWR _13381_ sky130_fd_sc_hd__mux2_1
X_22178_ _07361_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__buf_6
XFILLER_79_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21129_ _07776_ _07813_ _07814_ _07781_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__a22o_1
X_29774_ _13344_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__clkbuf_1
X_26986_ _11840_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__clkbuf_1
X_28725_ _12761_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__clkbuf_1
X_25937_ _11262_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28656_ _12725_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__clkbuf_1
X_16670_ _14998_ _15163_ _15166_ _15001_ VGND VGND VPWR VPWR _15167_ sky130_fd_sc_hd__a22o_1
X_25868_ _10858_ registers\[47\]\[61\] _11158_ VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__mux2_1
XFILLER_62_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27607_ registers\[34\]\[20\] _10346_ _12173_ VGND VGND VPWR VPWR _12174_ sky130_fd_sc_hd__mux2_1
X_24819_ _09613_ registers\[54\]\[47\] _10631_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__mux2_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28587_ _11807_ registers\[27\]\[37\] _12681_ VGND VGND VPWR VPWR _12689_ sky130_fd_sc_hd__mux2_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25799_ _10789_ registers\[47\]\[28\] _11181_ VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_404_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_404_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__buf_2
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27538_ _12136_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18271_ _14570_ _05033_ _05034_ _14582_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a22o_1
XFILLER_163_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ _12077_ VGND VGND VPWR VPWR _12100_ sky130_fd_sc_hd__buf_4
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29208_ registers\[23\]\[50\] _13039_ _13040_ VGND VGND VPWR VPWR _13041_ sky130_fd_sc_hd__mux2_1
XFILLER_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17222_ registers\[24\]\[32\] registers\[25\]\[32\] registers\[26\]\[32\] registers\[27\]\[32\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15704_ sky130_fd_sc_hd__mux4_1
XFILLER_230_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30480_ _13716_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 DW[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_6
Xinput25 DW[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
X_17153_ _15633_ _15634_ _15635_ _15636_ VGND VGND VPWR VPWR _15637_ sky130_fd_sc_hd__a22o_1
X_29139_ registers\[23\]\[28\] _12993_ _12977_ VGND VGND VPWR VPWR _12994_ sky130_fd_sc_hd__mux2_1
XFILLER_183_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 DW[41] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_4
XFILLER_156_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 DW[51] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_8
X_16104_ registers\[40\]\[1\] registers\[41\]\[1\] registers\[42\]\[1\] registers\[43\]\[1\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _14617_ sky130_fd_sc_hd__mux4_1
Xinput58 DW[61] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_16
Xinput69 R1[4] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
X_32150_ clknet_leaf_117_CLK _00264_ VGND VGND VPWR VPWR registers\[39\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_183_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17084_ _15295_ _15568_ _15569_ _15300_ VGND VGND VPWR VPWR _15570_ sky130_fd_sc_hd__a22o_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31101_ registers\[0\]\[45\] _13029_ _14037_ VGND VGND VPWR VPWR _14043_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16035_ _14548_ VGND VGND VPWR VPWR _14549_ sky130_fd_sc_hd__buf_4
X_32081_ clknet_leaf_491_CLK _00033_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31032_ registers\[0\]\[12\] _12960_ _14004_ VGND VGND VPWR VPWR _14007_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35840_ clknet_leaf_238_CLK _03954_ VGND VGND VPWR VPWR registers\[8\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_17986_ _04754_ _04758_ _04619_ _04620_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o211a_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19725_ _06374_ _06448_ _06449_ _06377_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__a22o_1
X_35771_ clknet_leaf_287_CLK _03885_ VGND VGND VPWR VPWR registers\[0\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_16937_ registers\[24\]\[24\] registers\[25\]\[24\] registers\[26\]\[24\] registers\[27\]\[24\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15427_ sky130_fd_sc_hd__mux4_1
X_32983_ clknet_leaf_62_CLK _01097_ VGND VGND VPWR VPWR registers\[52\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34722_ clknet_leaf_473_CLK _02836_ VGND VGND VPWR VPWR registers\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31934_ _09810_ registers\[49\]\[56\] _14474_ VGND VGND VPWR VPWR _14481_ sky130_fd_sc_hd__mux2_1
X_19656_ _06379_ _06380_ _06381_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__a22o_1
X_16868_ _15356_ _15359_ _15288_ VGND VGND VPWR VPWR _15360_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18607_ _05360_ _05363_ _05163_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__o21ba_1
XFILLER_80_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34653_ clknet_leaf_7_CLK _02767_ VGND VGND VPWR VPWR registers\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_19587_ _06312_ _06315_ _06180_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__o21ba_1
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31865_ _09730_ registers\[49\]\[23\] _14441_ VGND VGND VPWR VPWR _14445_ sky130_fd_sc_hd__mux2_1
X_16799_ _14597_ VGND VGND VPWR VPWR _15293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_241_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33604_ clknet_leaf_250_CLK _01718_ VGND VGND VPWR VPWR registers\[43\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_18538_ _05271_ _05280_ _05287_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__or4_4
X_30816_ _09771_ registers\[11\]\[38\] _13884_ VGND VGND VPWR VPWR _13893_ sky130_fd_sc_hd__mux2_1
XFILLER_244_1123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34584_ clknet_leaf_18_CLK _02698_ VGND VGND VPWR VPWR registers\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_31796_ _14408_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_233_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33535_ clknet_leaf_274_CLK _01649_ VGND VGND VPWR VPWR registers\[44\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18469_ registers\[20\]\[2\] registers\[21\]\[2\] registers\[22\]\[2\] registers\[23\]\[2\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30747_ _09668_ registers\[11\]\[5\] _13851_ VGND VGND VPWR VPWR _13857_ sky130_fd_sc_hd__mux2_1
XFILLER_142_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20500_ registers\[0\]\[61\] registers\[1\]\[61\] registers\[2\]\[61\] registers\[3\]\[61\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__mux4_1
XFILLER_222_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33466_ clknet_leaf_279_CLK _01580_ VGND VGND VPWR VPWR registers\[45\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21480_ registers\[40\]\[23\] registers\[41\]\[23\] registers\[42\]\[23\] registers\[43\]\[23\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__mux4_1
X_30678_ _13820_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35205_ clknet_leaf_220_CLK _03319_ VGND VGND VPWR VPWR registers\[18\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_20431_ _07131_ _07134_ _06847_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__o21ba_2
X_32417_ clknet_leaf_487_CLK _00531_ VGND VGND VPWR VPWR registers\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_36185_ clknet_leaf_92_CLK _00066_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33397_ clknet_leaf_344_CLK _01511_ VGND VGND VPWR VPWR registers\[46\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_35136_ clknet_leaf_240_CLK _03250_ VGND VGND VPWR VPWR registers\[1\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23150_ registers\[39\]\[20\] _09699_ _09700_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__mux2_1
X_20362_ _07065_ _07068_ _06880_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__o21ba_1
X_32348_ clknet_leaf_49_CLK _00462_ VGND VGND VPWR VPWR registers\[61\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22101_ _08755_ _08758_ _08759_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__o21ba_1
XTAP_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23081_ _09649_ _09650_ _09651_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__or3b_1
X_35067_ clknet_leaf_307_CLK _03181_ VGND VGND VPWR VPWR registers\[20\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_20293_ _06998_ _07001_ _06866_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__o21ba_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32279_ clknet_leaf_91_CLK _00393_ VGND VGND VPWR VPWR registers\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22032_ registers\[24\]\[38\] registers\[25\]\[38\] registers\[26\]\[38\] registers\[27\]\[38\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__mux4_1
X_34018_ clknet_leaf_48_CLK _02132_ VGND VGND VPWR VPWR registers\[36\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26840_ _11741_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_1
XTAP_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23983_ _09523_ registers\[5\]\[4\] _10161_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__mux2_1
X_26771_ _11657_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__buf_4
XFILLER_5_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35969_ clknet_leaf_231_CLK _04083_ VGND VGND VPWR VPWR registers\[6\]\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_229_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28510_ _11728_ registers\[27\]\[0\] _12648_ VGND VGND VPWR VPWR _12649_ sky130_fd_sc_hd__mux2_1
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25722_ _11148_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22934_ _09551_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
X_29490_ _13139_ VGND VGND VPWR VPWR _13195_ sky130_fd_sc_hd__buf_4
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28441_ _12612_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__clkbuf_1
X_22865_ _09497_ _09500_ _07369_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__o21ba_1
XFILLER_3_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25653_ _11112_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21816_ registers\[0\]\[32\] registers\[1\]\[32\] registers\[2\]\[32\] registers\[3\]\[32\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__mux4_1
X_24604_ _10513_ VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__clkbuf_8
X_28372_ _12575_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__clkbuf_1
X_25584_ _11074_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22796_ registers\[52\]\[61\] registers\[53\]\[61\] registers\[54\]\[61\] registers\[55\]\[61\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__mux4_1
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_974 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24535_ _10487_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
X_27323_ _12023_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__clkbuf_1
X_21747_ _07369_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__clkbuf_4
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27254_ _11826_ registers\[37\]\[46\] _11980_ VGND VGND VPWR VPWR _11987_ sky130_fd_sc_hd__mux2_1
X_24466_ _10439_ VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__buf_4
XFILLER_196_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21678_ _08343_ _08348_ _08073_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__o21ba_1
XFILLER_40_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23417_ registers\[39\]\[61\] _09821_ _09657_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__mux2_1
X_26205_ _11403_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
X_20629_ _07280_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__buf_12
X_27185_ _11757_ registers\[37\]\[13\] _11947_ VGND VGND VPWR VPWR _11951_ sky130_fd_sc_hd__mux2_1
X_24397_ net44 VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__buf_4
XFILLER_138_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26136_ _10856_ registers\[45\]\[60\] _11300_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__mux2_1
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23348_ registers\[39\]\[28\] _09749_ _09700_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26067_ _10787_ registers\[45\]\[27\] _11323_ VGND VGND VPWR VPWR _11331_ sky130_fd_sc_hd__mux2_1
XFILLER_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23279_ _09781_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_1
X_25018_ _10748_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1604 _14567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1615 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1626 _15845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17840_ registers\[52\]\[50\] registers\[53\]\[50\] registers\[54\]\[50\] registers\[55\]\[50\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__mux4_1
XFILLER_152_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1637 net260 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29826_ registers\[18\]\[17\] _12970_ _13364_ VGND VGND VPWR VPWR _13372_ sky130_fd_sc_hd__mux2_1
XTAP_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1648 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1659 _00028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17771_ registers\[60\]\[48\] registers\[61\]\[48\] registers\[62\]\[48\] registers\[63\]\[48\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__mux4_1
X_29757_ _13335_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__clkbuf_1
X_26969_ _11828_ registers\[3\]\[47\] _11814_ VGND VGND VPWR VPWR _11829_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_1375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19510_ _06090_ _06239_ _06240_ _06096_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__a22o_1
XFILLER_47_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16722_ _14578_ VGND VGND VPWR VPWR _15218_ sky130_fd_sc_hd__buf_4
X_28708_ _11792_ registers\[26\]\[30\] _12752_ VGND VGND VPWR VPWR _12753_ sky130_fd_sc_hd__mux2_1
XFILLER_235_633 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29688_ _13299_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19441_ _05113_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__buf_4
X_28639_ _11859_ registers\[27\]\[62\] _12647_ VGND VGND VPWR VPWR _12716_ sky130_fd_sc_hd__mux2_1
XFILLER_223_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16653_ _14592_ VGND VGND VPWR VPWR _15151_ sky130_fd_sc_hd__buf_6
XFILLER_228_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_1419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31650_ _14331_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__clkbuf_1
X_19372_ _06031_ _06105_ _06106_ _06034_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__a22o_1
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16584_ registers\[24\]\[14\] registers\[25\]\[14\] registers\[26\]\[14\] registers\[27\]\[14\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15084_ sky130_fd_sc_hd__mux4_1
XFILLER_215_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18323_ _05049_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__buf_2
X_30601_ _13779_ VGND VGND VPWR VPWR _13780_ sky130_fd_sc_hd__buf_4
XFILLER_128_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31581_ _14295_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__clkbuf_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_787 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33320_ clknet_leaf_59_CLK _01434_ VGND VGND VPWR VPWR registers\[47\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18254_ _14587_ _05016_ _05017_ _14597_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__a22o_1
X_30532_ _09756_ registers\[13\]\[31\] _13742_ VGND VGND VPWR VPWR _13744_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17205_ _14516_ VGND VGND VPWR VPWR _15687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33251_ clknet_leaf_47_CLK _01365_ VGND VGND VPWR VPWR registers\[48\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_30463_ _09825_ registers\[14\]\[63\] _13637_ VGND VGND VPWR VPWR _13707_ sky130_fd_sc_hd__mux2_1
X_18185_ registers\[40\]\[61\] registers\[41\]\[61\] registers\[42\]\[61\] registers\[43\]\[61\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__mux4_1
XFILLER_204_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32202_ clknet_leaf_380_CLK _00316_ VGND VGND VPWR VPWR registers\[9\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17136_ _14553_ VGND VGND VPWR VPWR _15620_ sky130_fd_sc_hd__clkbuf_4
X_33182_ clknet_leaf_477_CLK _01296_ VGND VGND VPWR VPWR registers\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30394_ _13637_ VGND VGND VPWR VPWR _13671_ sky130_fd_sc_hd__buf_6
XFILLER_183_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32133_ clknet_leaf_460_CLK _00050_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17067_ _14516_ VGND VGND VPWR VPWR _15553_ sky130_fd_sc_hd__clkbuf_8
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16018_ _14531_ VGND VGND VPWR VPWR _14532_ sky130_fd_sc_hd__buf_4
X_32064_ clknet_leaf_294_CLK _00242_ VGND VGND VPWR VPWR registers\[62\]\[50\] sky130_fd_sc_hd__dfxtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_890 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31015_ registers\[0\]\[4\] _12943_ _13993_ VGND VGND VPWR VPWR _13998_ sky130_fd_sc_hd__mux2_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35823_ clknet_leaf_376_CLK _03937_ VGND VGND VPWR VPWR registers\[8\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_17969_ _04719_ _04726_ _04735_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__or4_4
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19708_ _05076_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__clkbuf_4
X_35754_ clknet_leaf_399_CLK _03868_ VGND VGND VPWR VPWR registers\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_32966_ clknet_leaf_194_CLK _01080_ VGND VGND VPWR VPWR registers\[53\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20980_ _07639_ _07654_ _07663_ _07670_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__or4_1
XFILLER_84_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34705_ clknet_leaf_111_CLK _02819_ VGND VGND VPWR VPWR registers\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31917_ _09793_ registers\[49\]\[48\] _14463_ VGND VGND VPWR VPWR _14472_ sky130_fd_sc_hd__mux2_1
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19639_ registers\[48\]\[36\] registers\[49\]\[36\] registers\[50\]\[36\] registers\[51\]\[36\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux4_1
Xclkbuf_2_2_0_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_2_0_CLK sky130_fd_sc_hd__clkbuf_8
X_35685_ clknet_leaf_465_CLK _03799_ VGND VGND VPWR VPWR registers\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_32897_ clknet_leaf_294_CLK _01011_ VGND VGND VPWR VPWR registers\[54\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34636_ clknet_leaf_148_CLK _02750_ VGND VGND VPWR VPWR registers\[27\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_22650_ registers\[0\]\[56\] registers\[1\]\[56\] registers\[2\]\[56\] registers\[3\]\[56\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1027 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31848_ _09689_ registers\[49\]\[15\] _14430_ VGND VGND VPWR VPWR _14436_ sky130_fd_sc_hd__mux2_1
X_21601_ registers\[4\]\[26\] registers\[5\]\[26\] registers\[6\]\[26\] registers\[7\]\[26\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__mux4_1
XFILLER_209_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34567_ clknet_leaf_206_CLK _02681_ VGND VGND VPWR VPWR registers\[28\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_22581_ _09012_ _09224_ _09225_ _09018_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__a22o_1
XFILLER_90_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31779_ _14399_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24320_ net17 VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__clkbuf_4
X_21532_ registers\[4\]\[24\] registers\[5\]\[24\] registers\[6\]\[24\] registers\[7\]\[24\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__mux4_1
X_33518_ clknet_leaf_361_CLK _01632_ VGND VGND VPWR VPWR registers\[44\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34498_ clknet_leaf_241_CLK _02612_ VGND VGND VPWR VPWR registers\[2\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36237_ clknet_leaf_122_CLK _00123_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dfxtp_1
X_24251_ _10308_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
X_33449_ clknet_leaf_60_CLK _01563_ VGND VGND VPWR VPWR registers\[45\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_21463_ registers\[0\]\[22\] registers\[1\]\[22\] registers\[2\]\[22\] registers\[3\]\[22\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__mux4_1
X_23202_ registers\[9\]\[17\] _09693_ _09722_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__mux2_1
X_20414_ _05060_ _07117_ _07118_ _05066_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36168_ clknet_leaf_193_CLK _04282_ VGND VGND VPWR VPWR registers\[49\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_24182_ _09586_ registers\[58\]\[34\] _10266_ VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__mux2_1
XFILLER_175_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21394_ _07369_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__buf_2
XFILLER_147_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35119_ clknet_leaf_377_CLK _03233_ VGND VGND VPWR VPWR registers\[1\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_23133_ net7 VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__buf_6
X_20345_ registers\[60\]\[56\] registers\[61\]\[56\] registers\[62\]\[56\] registers\[63\]\[56\]
+ _06991_ _06785_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__mux4_1
X_36099_ clknet_leaf_263_CLK _04213_ VGND VGND VPWR VPWR registers\[59\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28990_ registers\[24\]\[36\] _10380_ _12894_ VGND VGND VPWR VPWR _12901_ sky130_fd_sc_hd__mux2_1
XFILLER_162_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27941_ _12349_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__clkbuf_1
X_23064_ _09639_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20276_ _06919_ _06983_ _06984_ _06922_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__a22o_1
XTAP_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22015_ _08669_ _08671_ _08674_ _08675_ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__a22o_1
XTAP_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27872_ registers\[32\]\[18\] _10342_ _12304_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__mux2_1
XTAP_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29611_ registers\[20\]\[43\] _13025_ _13255_ VGND VGND VPWR VPWR _13259_ sky130_fd_sc_hd__mux2_1
XFILLER_248_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _11729_ VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__buf_4
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29542_ registers\[20\]\[10\] _12955_ _13222_ VGND VGND VPWR VPWR _13223_ sky130_fd_sc_hd__mux2_1
XFILLER_229_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26754_ _11693_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_1
X_23966_ _09642_ registers\[60\]\[61\] _10088_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__mux2_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25705_ _11139_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
X_29473_ _13186_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__clkbuf_1
X_22917_ net4 VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__buf_4
X_26685_ _11084_ _11157_ VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__and2b_1
XFILLER_217_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23897_ _09573_ registers\[60\]\[28\] _10111_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__mux2_1
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28424_ _12603_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__clkbuf_1
X_22848_ registers\[44\]\[63\] registers\[45\]\[63\] registers\[46\]\[63\] registers\[47\]\[63\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__mux4_1
X_25636_ _11103_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28355_ registers\[2\]\[55\] _10420_ _12561_ VGND VGND VPWR VPWR _12567_ sky130_fd_sc_hd__mux2_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ registers\[28\]\[60\] registers\[29\]\[60\] registers\[30\]\[60\] registers\[31\]\[60\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__mux4_1
XFILLER_197_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25567_ _11065_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27306_ _12014_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24518_ _10478_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28286_ registers\[2\]\[22\] _10351_ _12528_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__mux2_1
X_25498_ _11029_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_1
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27237_ _11809_ registers\[37\]\[38\] _11969_ VGND VGND VPWR VPWR _11978_ sky130_fd_sc_hd__mux2_1
X_24449_ _10442_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27168_ _11740_ registers\[37\]\[5\] _11936_ VGND VGND VPWR VPWR _11942_ sky130_fd_sc_hd__mux2_1
XFILLER_165_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26119_ _11358_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
X_19990_ _06703_ _06706_ _06504_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__o21ba_1
XFILLER_126_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27099_ _11905_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18941_ _05039_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1401 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1412 _00179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1423 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18872_ registers\[52\]\[14\] registers\[53\]\[14\] registers\[54\]\[14\] registers\[55\]\[14\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__mux4_1
XFILLER_45_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1434 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1445 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1456 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17823_ _04597_ _04600_ _04301_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29809_ registers\[18\]\[9\] _12953_ _13353_ VGND VGND VPWR VPWR _13363_ sky130_fd_sc_hd__mux2_1
XTAP_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1467 _05162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1478 _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1489 _07309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32820_ clknet_leaf_352_CLK _00934_ VGND VGND VPWR VPWR registers\[55\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17754_ registers\[40\]\[48\] registers\[41\]\[48\] registers\[42\]\[48\] registers\[43\]\[48\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__mux4_1
XTAP_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16705_ _14493_ VGND VGND VPWR VPWR _15201_ sky130_fd_sc_hd__buf_4
X_32751_ clknet_leaf_367_CLK _00865_ VGND VGND VPWR VPWR registers\[56\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17685_ registers\[32\]\[46\] registers\[33\]\[46\] registers\[34\]\[46\] registers\[35\]\[46\]
+ _15917_ _15918_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__mux4_1
XFILLER_90_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19424_ _05097_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__clkbuf_4
X_31702_ _14347_ VGND VGND VPWR VPWR _14359_ sky130_fd_sc_hd__buf_4
X_35470_ clknet_leaf_137_CLK _03584_ VGND VGND VPWR VPWR registers\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16636_ _14546_ VGND VGND VPWR VPWR _15134_ sky130_fd_sc_hd__clkbuf_8
X_32682_ clknet_leaf_424_CLK _00796_ VGND VGND VPWR VPWR registers\[57\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34421_ clknet_leaf_416_CLK _02535_ VGND VGND VPWR VPWR registers\[30\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_19355_ _05076_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__buf_4
XFILLER_91_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31633_ registers\[63\]\[41\] net36 _14321_ VGND VGND VPWR VPWR _14323_ sky130_fd_sc_hd__mux2_1
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16567_ registers\[56\]\[14\] registers\[57\]\[14\] registers\[58\]\[14\] registers\[59\]\[14\]
+ _15066_ _14856_ VGND VGND VPWR VPWR _15067_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18306_ _05044_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__buf_12
X_34352_ clknet_leaf_387_CLK _02466_ VGND VGND VPWR VPWR registers\[31\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31564_ _14286_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19286_ registers\[48\]\[26\] registers\[49\]\[26\] registers\[50\]\[26\] registers\[51\]\[26\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__mux4_1
XFILLER_175_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16498_ registers\[36\]\[12\] registers\[37\]\[12\] registers\[38\]\[12\] registers\[39\]\[12\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _15000_ sky130_fd_sc_hd__mux4_1
XFILLER_148_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33303_ clknet_leaf_123_CLK _01417_ VGND VGND VPWR VPWR registers\[47\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18237_ registers\[16\]\[62\] registers\[17\]\[62\] registers\[18\]\[62\] registers\[19\]\[62\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__mux4_1
X_30515_ _09730_ registers\[13\]\[23\] _13731_ VGND VGND VPWR VPWR _13735_ sky130_fd_sc_hd__mux2_1
X_34283_ clknet_leaf_426_CLK _02397_ VGND VGND VPWR VPWR registers\[32\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_31495_ _14205_ VGND VGND VPWR VPWR _14250_ sky130_fd_sc_hd__buf_4
XFILLER_50_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36022_ clknet_leaf_330_CLK _04136_ VGND VGND VPWR VPWR registers\[63\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33234_ clknet_leaf_74_CLK _01348_ VGND VGND VPWR VPWR registers\[48\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30446_ _13698_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__clkbuf_1
X_18168_ _04931_ _04934_ _14553_ _14555_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__o211a_1
XFILLER_175_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17119_ _15603_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
X_33165_ clknet_leaf_170_CLK _01279_ VGND VGND VPWR VPWR registers\[50\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18099_ registers\[36\]\[58\] registers\[37\]\[58\] registers\[38\]\[58\] registers\[39\]\[58\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__mux4_1
XFILLER_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30377_ _13662_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__clkbuf_1
X_20130_ _05097_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32116_ clknet_leaf_467_CLK _00031_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dfxtp_1
X_33096_ clknet_leaf_194_CLK _01210_ VGND VGND VPWR VPWR registers\[51\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20061_ _05038_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__clkbuf_4
X_32047_ clknet_leaf_370_CLK _00225_ VGND VGND VPWR VPWR registers\[62\]\[33\] sky130_fd_sc_hd__dfxtp_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23820_ _09632_ registers\[29\]\[56\] _10072_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__mux2_1
XFILLER_113_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35806_ clknet_leaf_485_CLK _03920_ VGND VGND VPWR VPWR registers\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33998_ clknet_leaf_133_CLK _02112_ VGND VGND VPWR VPWR registers\[36\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _09563_ registers\[29\]\[23\] _10039_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__mux2_1
X_20963_ _07647_ _07653_ _07339_ _07341_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__o211a_1
XANTENNA_309 _00087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35737_ clknet_leaf_13_CLK _03851_ VGND VGND VPWR VPWR registers\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_32949_ clknet_leaf_352_CLK _01063_ VGND VGND VPWR VPWR registers\[53\]\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22702_ registers\[56\]\[58\] registers\[57\]\[58\] registers\[58\]\[58\] registers\[59\]\[58\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__mux4_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23682_ registers\[61\]\[56\] _09810_ _09998_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__mux2_1
X_26470_ _10785_ registers\[42\]\[26\] _11536_ VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__mux2_1
X_20894_ registers\[12\]\[6\] registers\[13\]\[6\] registers\[14\]\[6\] registers\[15\]\[6\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__mux4_1
X_35668_ clknet_leaf_88_CLK _03782_ VGND VGND VPWR VPWR registers\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22633_ _09255_ _09262_ _09269_ _09276_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__or4_4
X_25421_ _10825_ registers\[50\]\[45\] _10981_ VGND VGND VPWR VPWR _10987_ sky130_fd_sc_hd__mux2_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34619_ clknet_leaf_183_CLK _02733_ VGND VGND VPWR VPWR registers\[27\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35599_ clknet_leaf_134_CLK _03713_ VGND VGND VPWR VPWR registers\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25352_ _10756_ registers\[50\]\[12\] _10948_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__mux2_1
X_28140_ _11765_ registers\[30\]\[17\] _12446_ VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__mux2_1
X_22564_ _09104_ _09208_ _09209_ _09107_ VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__a22o_1
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21515_ registers\[44\]\[24\] registers\[45\]\[24\] registers\[46\]\[24\] registers\[47\]\[24\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__mux4_1
XFILLER_22_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24303_ _10343_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
X_28071_ _12417_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__clkbuf_1
X_25283_ _10823_ registers\[51\]\[44\] _10909_ VGND VGND VPWR VPWR _10914_ sky130_fd_sc_hd__mux2_1
XFILLER_107_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22495_ registers\[28\]\[51\] registers\[29\]\[51\] registers\[30\]\[51\] registers\[31\]\[51\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27022_ _11864_ VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__buf_4
X_24234_ _09638_ registers\[58\]\[59\] _10288_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__mux2_1
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21446_ registers\[32\]\[22\] registers\[33\]\[22\] registers\[34\]\[22\] registers\[35\]\[22\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__mux4_1
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24165_ _09569_ registers\[58\]\[26\] _10255_ VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__mux2_1
XFILLER_218_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21377_ registers\[56\]\[20\] registers\[57\]\[20\] registers\[58\]\[20\] registers\[59\]\[20\]
+ _07851_ _07984_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__mux4_1
XFILLER_218_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23116_ _09677_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
X_20328_ _06868_ _07034_ _07035_ _06871_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__a22o_1
XFILLER_150_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24096_ _09636_ registers\[5\]\[58\] _10216_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__mux2_1
X_28973_ registers\[24\]\[28\] _10363_ _12883_ VGND VGND VPWR VPWR _12892_ sky130_fd_sc_hd__mux2_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23047_ net50 VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__buf_4
X_27924_ _12340_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_1
X_20259_ registers\[4\]\[53\] registers\[5\]\[53\] registers\[6\]\[53\] registers\[7\]\[53\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux4_1
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27855_ _12292_ VGND VGND VPWR VPWR _12304_ sky130_fd_sc_hd__buf_6
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_1__f_CLK clknet_5_0_0_CLK VGND VGND VPWR VPWR clknet_6_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26806_ _11720_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__clkbuf_1
XTAP_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27786_ registers\[33\]\[41\] _10391_ _12266_ VGND VGND VPWR VPWR _12268_ sky130_fd_sc_hd__mux2_1
X_24998_ net23 VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__buf_4
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29525_ registers\[20\]\[2\] _12939_ _13211_ VGND VGND VPWR VPWR _13214_ sky130_fd_sc_hd__mux2_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26737_ _11684_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__clkbuf_1
X_23949_ _10147_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_245_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_810 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_821 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_832 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29456_ _13177_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__clkbuf_1
X_17470_ _15941_ _15944_ _15645_ VGND VGND VPWR VPWR _15945_ sky130_fd_sc_hd__o21ba_1
X_26668_ _11647_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_843 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_854 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_865 _09335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_232_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16421_ _14655_ _14923_ _14924_ _14658_ VGND VGND VPWR VPWR _14925_ sky130_fd_sc_hd__a22o_1
X_28407_ _12594_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25619_ _11094_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_876 _09527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_847 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29387_ _13141_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_887 _09611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_898 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26599_ _11611_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19140_ _05860_ _05867_ _05874_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__or4_2
X_28338_ registers\[2\]\[47\] _10403_ _12550_ VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__mux2_1
X_16352_ _14493_ VGND VGND VPWR VPWR _14858_ sky130_fd_sc_hd__buf_4
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19071_ _05097_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__clkbuf_4
X_16283_ _14546_ VGND VGND VPWR VPWR _14791_ sky130_fd_sc_hd__buf_4
XFILLER_9_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28269_ registers\[2\]\[14\] _10334_ _12517_ VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__mux2_1
XFILLER_200_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30300_ _13565_ VGND VGND VPWR VPWR _13621_ sky130_fd_sc_hd__buf_4
X_18022_ registers\[12\]\[55\] registers\[13\]\[55\] registers\[14\]\[55\] registers\[15\]\[55\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux4_1
XFILLER_172_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31280_ _14137_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_952 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30231_ registers\[15\]\[17\] _12970_ _13577_ VGND VGND VPWR VPWR _13585_ sky130_fd_sc_hd__mux2_1
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30162_ _13548_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__clkbuf_1
X_19973_ _06379_ _06689_ _06690_ _06382_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__a22o_1
XFILLER_10_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18924_ _05671_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34970_ clknet_leaf_0_CLK _03084_ VGND VGND VPWR VPWR registers\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1220 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30093_ _13512_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1231 _00034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1242 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33921_ clknet_leaf_258_CLK _02035_ VGND VGND VPWR VPWR registers\[38\]\[51\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1253 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18855_ _05501_ _05603_ _05604_ _05506_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__a22o_1
XTAP_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1264 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1275 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1286 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ registers\[60\]\[49\] registers\[61\]\[49\] registers\[62\]\[49\] registers\[63\]\[49\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__mux4_1
XFILLER_83_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1297 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33852_ clknet_leaf_299_CLK _01966_ VGND VGND VPWR VPWR registers\[3\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18786_ _05534_ _05537_ _05508_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__o21ba_1
X_15998_ _14502_ VGND VGND VPWR VPWR _14512_ sky130_fd_sc_hd__buf_4
XTAP_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32803_ clknet_leaf_443_CLK _00917_ VGND VGND VPWR VPWR registers\[55\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17737_ _04513_ _04516_ _15963_ _15964_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__o211a_1
XFILLER_76_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33783_ clknet_leaf_341_CLK _01897_ VGND VGND VPWR VPWR registers\[40\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_30995_ registers\[10\]\[59\] _13058_ _13977_ VGND VGND VPWR VPWR _13987_ sky130_fd_sc_hd__mux2_1
XFILLER_223_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35522_ clknet_leaf_238_CLK _03636_ VGND VGND VPWR VPWR registers\[13\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32734_ clknet_leaf_38_CLK _00848_ VGND VGND VPWR VPWR registers\[56\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_17668_ registers\[8\]\[45\] registers\[9\]\[45\] registers\[10\]\[45\] registers\[11\]\[45\]
+ _04448_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__mux4_1
XFILLER_247_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19407_ registers\[12\]\[29\] registers\[13\]\[29\] registers\[14\]\[29\] registers\[15\]\[29\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__mux4_1
X_35453_ clknet_leaf_298_CLK _03567_ VGND VGND VPWR VPWR registers\[14\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_16619_ registers\[28\]\[15\] registers\[29\]\[15\] registers\[30\]\[15\] registers\[31\]\[15\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15118_ sky130_fd_sc_hd__mux4_1
X_32665_ clknet_leaf_84_CLK _00779_ VGND VGND VPWR VPWR registers\[57\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17599_ _04379_ _04382_ _15963_ _15964_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__o211a_1
XFILLER_204_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34404_ clknet_leaf_472_CLK _02518_ VGND VGND VPWR VPWR registers\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_19338_ _06070_ _06073_ _05837_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__o21ba_1
X_31616_ registers\[63\]\[33\] net27 _14310_ VGND VGND VPWR VPWR _14314_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35384_ clknet_leaf_320_CLK _03498_ VGND VGND VPWR VPWR registers\[15\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32596_ clknet_leaf_71_CLK _00710_ VGND VGND VPWR VPWR registers\[58\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_34335_ clknet_leaf_488_CLK _02449_ VGND VGND VPWR VPWR registers\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31547_ registers\[63\]\[0\] net1 _14277_ VGND VGND VPWR VPWR _14278_ sky130_fd_sc_hd__mux2_1
XFILLER_149_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19269_ registers\[24\]\[25\] registers\[25\]\[25\] registers\[26\]\[25\] registers\[27\]\[25\]
+ _05974_ _05975_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__mux4_1
XFILLER_143_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21300_ _07783_ _07979_ _07980_ _07786_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__a22o_1
XFILLER_178_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22280_ _08766_ _08932_ _08933_ _08771_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__a22o_1
X_34266_ clknet_leaf_18_CLK _02380_ VGND VGND VPWR VPWR registers\[32\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_31478_ _14241_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__clkbuf_1
X_36005_ clknet_leaf_450_CLK _04119_ VGND VGND VPWR VPWR registers\[63\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_33217_ clknet_leaf_234_CLK _01331_ VGND VGND VPWR VPWR registers\[4\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_21231_ _07910_ _07913_ _07711_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__o21ba_1
XFILLER_176_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30429_ _13689_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__clkbuf_1
X_34197_ clknet_leaf_122_CLK _02311_ VGND VGND VPWR VPWR registers\[33\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33148_ clknet_leaf_276_CLK _01262_ VGND VGND VPWR VPWR registers\[50\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_21162_ registers\[44\]\[14\] registers\[45\]\[14\] registers\[46\]\[14\] registers\[47\]\[14\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__mux4_1
XFILLER_105_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20113_ registers\[12\]\[49\] registers\[13\]\[49\] registers\[14\]\[49\] registers\[15\]\[49\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__mux4_1
XFILLER_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25970_ _10825_ registers\[46\]\[45\] _11274_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__mux2_1
X_21093_ registers\[32\]\[12\] registers\[33\]\[12\] registers\[34\]\[12\] registers\[35\]\[12\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__mux4_1
X_33079_ clknet_leaf_343_CLK _01193_ VGND VGND VPWR VPWR registers\[51\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_217_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20044_ _06756_ _06759_ _06523_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__o21ba_1
X_24921_ _09580_ registers\[53\]\[31\] _10691_ VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__mux2_1
XFILLER_219_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_213_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27640_ registers\[34\]\[36\] _10380_ _12184_ VGND VGND VPWR VPWR _12191_ sky130_fd_sc_hd__mux2_1
XFILLER_100_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24852_ _09646_ registers\[54\]\[63\] _10586_ VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__mux2_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23803_ _09615_ registers\[29\]\[48\] _10061_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__mux2_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27571_ registers\[34\]\[3\] _10311_ _12151_ VGND VGND VPWR VPWR _12155_ sky130_fd_sc_hd__mux2_1
XFILLER_233_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ registers\[28\]\[37\] registers\[29\]\[37\] registers\[30\]\[37\] registers\[31\]\[37\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__mux4_1
X_24783_ _10586_ VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__clkbuf_8
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_117 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29310_ _13100_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26522_ _11570_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_128 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ registers\[36\]\[8\] registers\[37\]\[8\] registers\[38\]\[8\] registers\[39\]\[8\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__mux4_1
X_23734_ _09546_ registers\[29\]\[15\] _10028_ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__mux2_1
XANTENNA_139 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29241_ registers\[23\]\[61\] _13062_ _12934_ VGND VGND VPWR VPWR _13063_ sky130_fd_sc_hd__mux2_1
XFILLER_121_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26453_ _10768_ registers\[42\]\[18\] _11525_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__mux2_1
X_20877_ _07440_ _07568_ _07569_ _07443_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__a22o_1
X_23665_ registers\[61\]\[48\] _09793_ _09987_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__mux2_1
XFILLER_14_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25404_ _10808_ registers\[50\]\[37\] _10970_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__mux2_1
X_22616_ registers\[52\]\[55\] registers\[53\]\[55\] registers\[54\]\[55\] registers\[55\]\[55\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__mux4_1
X_29172_ net33 VGND VGND VPWR VPWR _13016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26384_ _11497_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__clkbuf_1
X_23596_ registers\[61\]\[15\] _09689_ _09954_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__mux2_1
XFILLER_167_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28123_ _11748_ registers\[30\]\[9\] _12435_ VGND VGND VPWR VPWR _12445_ sky130_fd_sc_hd__mux2_1
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22547_ registers\[48\]\[53\] registers\[49\]\[53\] registers\[50\]\[53\] registers\[51\]\[53\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__mux4_1
X_25335_ _10739_ registers\[50\]\[4\] _10937_ VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__mux2_1
XFILLER_128_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28054_ _11813_ registers\[31\]\[40\] _12408_ VGND VGND VPWR VPWR _12409_ sky130_fd_sc_hd__mux2_1
X_22478_ registers\[56\]\[51\] registers\[57\]\[51\] registers\[58\]\[51\] registers\[59\]\[51\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__mux4_1
XFILLER_155_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25266_ _10806_ registers\[51\]\[36\] _10898_ VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__mux2_1
XFILLER_136_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27005_ net55 VGND VGND VPWR VPWR _11853_ sky130_fd_sc_hd__clkbuf_4
X_24217_ _10289_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
X_21429_ registers\[12\]\[21\] registers\[13\]\[21\] registers\[14\]\[21\] registers\[15\]\[21\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__mux4_1
X_25197_ _10737_ registers\[51\]\[3\] _10865_ VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__mux2_1
XFILLER_163_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_922 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24148_ _09552_ registers\[58\]\[18\] _10244_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__mux2_1
XFILLER_159_1384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24079_ _10160_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__buf_4
X_16970_ registers\[16\]\[25\] registers\[17\]\[25\] registers\[18\]\[25\] registers\[19\]\[25\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15459_ sky130_fd_sc_hd__mux4_1
X_28956_ net282 VGND VGND VPWR VPWR _12883_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27907_ _12331_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__clkbuf_1
X_28887_ _11837_ registers\[25\]\[51\] _12845_ VGND VGND VPWR VPWR _12847_ sky130_fd_sc_hd__mux2_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _05374_ _05381_ _05388_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__or4_4
X_27838_ _12295_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__clkbuf_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _05328_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27769_ registers\[33\]\[33\] _10374_ _12255_ VGND VGND VPWR VPWR _12259_ sky130_fd_sc_hd__mux2_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29508_ _13204_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__clkbuf_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ registers\[36\]\[41\] registers\[37\]\[41\] registers\[38\]\[41\] registers\[39\]\[41\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__mux4_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30780_ _13874_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__clkbuf_1
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_640 _05156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_651 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_662 _05297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29439_ _13168_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__clkbuf_1
X_17453_ registers\[60\]\[39\] registers\[61\]\[39\] registers\[62\]\[39\] registers\[63\]\[39\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _15928_ sky130_fd_sc_hd__mux4_1
XANTENNA_673 _05687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_684 _06195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_695 _07135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16404_ _14905_ _14908_ _14585_ VGND VGND VPWR VPWR _14909_ sky130_fd_sc_hd__o21ba_1
X_32450_ clknet_leaf_229_CLK _00564_ VGND VGND VPWR VPWR registers\[29\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_17384_ _15857_ _15860_ _15620_ _15621_ VGND VGND VPWR VPWR _15861_ sky130_fd_sc_hd__o211a_1
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31401_ _14200_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__clkbuf_1
X_19123_ registers\[52\]\[21\] registers\[53\]\[21\] registers\[54\]\[21\] registers\[55\]\[21\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__mux4_1
X_16335_ _14588_ _14840_ _14841_ _14598_ VGND VGND VPWR VPWR _14842_ sky130_fd_sc_hd__a22o_1
XFILLER_207_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32381_ clknet_leaf_288_CLK _00495_ VGND VGND VPWR VPWR registers\[61\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34120_ clknet_leaf_244_CLK _02234_ VGND VGND VPWR VPWR registers\[35\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31332_ _14164_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__clkbuf_1
X_19054_ registers\[12\]\[19\] registers\[13\]\[19\] registers\[14\]\[19\] registers\[15\]\[19\]
+ _05594_ _05595_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__mux4_1
X_16266_ registers\[28\]\[5\] registers\[29\]\[5\] registers\[30\]\[5\] registers\[31\]\[5\]
+ _14678_ _14679_ VGND VGND VPWR VPWR _14775_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18005_ registers\[40\]\[55\] registers\[41\]\[55\] registers\[42\]\[55\] registers\[43\]\[55\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__mux4_1
X_34051_ clknet_leaf_251_CLK _02165_ VGND VGND VPWR VPWR registers\[36\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_31263_ registers\[8\]\[58\] net54 _14119_ VGND VGND VPWR VPWR _14128_ sky130_fd_sc_hd__mux2_1
X_16197_ registers\[24\]\[3\] registers\[25\]\[3\] registers\[26\]\[3\] registers\[27\]\[3\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _14708_ sky130_fd_sc_hd__mux4_1
XFILLER_12_1277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33002_ clknet_leaf_422_CLK _01116_ VGND VGND VPWR VPWR registers\[52\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30214_ registers\[15\]\[9\] _12953_ _13566_ VGND VGND VPWR VPWR _13576_ sky130_fd_sc_hd__mux2_1
XFILLER_126_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31194_ registers\[8\]\[25\] net18 _14086_ VGND VGND VPWR VPWR _14092_ sky130_fd_sc_hd__mux2_1
XFILLER_181_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30145_ registers\[16\]\[40\] _13018_ _13539_ VGND VGND VPWR VPWR _13540_ sky130_fd_sc_hd__mux2_1
X_19956_ registers\[36\]\[45\] registers\[37\]\[45\] registers\[38\]\[45\] registers\[39\]\[45\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__mux4_1
XFILLER_114_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18907_ _05051_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__buf_4
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34953_ clknet_leaf_212_CLK _03067_ VGND VGND VPWR VPWR registers\[22\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_30076_ _13503_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1050 _13423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19887_ registers\[32\]\[43\] registers\[33\]\[43\] registers\[34\]\[43\] registers\[35\]\[43\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__mux4_1
XFILLER_206_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1061 _13992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_210_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1072 _14347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1083 _14499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33904_ clknet_leaf_357_CLK _02018_ VGND VGND VPWR VPWR registers\[38\]\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1094 _14524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18838_ registers\[52\]\[13\] registers\[53\]\[13\] registers\[54\]\[13\] registers\[55\]\[13\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__mux4_1
XFILLER_3_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34884_ clknet_leaf_203_CLK _02998_ VGND VGND VPWR VPWR registers\[23\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18769_ registers\[60\]\[11\] registers\[61\]\[11\] registers\[62\]\[11\] registers\[63\]\[11\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__mux4_1
X_33835_ clknet_leaf_458_CLK _01949_ VGND VGND VPWR VPWR registers\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20800_ registers\[28\]\[3\] registers\[29\]\[3\] registers\[30\]\[3\] registers\[31\]\[3\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__mux4_1
XFILLER_82_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21780_ registers\[0\]\[31\] registers\[1\]\[31\] registers\[2\]\[31\] registers\[3\]\[31\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__mux4_1
X_33766_ clknet_leaf_432_CLK _01880_ VGND VGND VPWR VPWR registers\[40\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_30978_ _13978_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20731_ registers\[20\]\[1\] registers\[21\]\[1\] registers\[22\]\[1\] registers\[23\]\[1\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__mux4_1
XFILLER_19_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35505_ clknet_leaf_378_CLK _03619_ VGND VGND VPWR VPWR registers\[13\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32717_ clknet_leaf_139_CLK _00831_ VGND VGND VPWR VPWR registers\[57\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33697_ clknet_leaf_39_CLK _01811_ VGND VGND VPWR VPWR registers\[41\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23450_ _09882_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__clkbuf_1
X_32648_ clknet_leaf_209_CLK _00762_ VGND VGND VPWR VPWR registers\[58\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_35436_ clknet_leaf_394_CLK _03550_ VGND VGND VPWR VPWR registers\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_20662_ _07314_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__buf_12
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22401_ _08812_ _09049_ _09050_ _08815_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__a22o_1
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23381_ _09844_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
X_20593_ _07276_ _07283_ _07286_ _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__a22o_1
X_32579_ clknet_leaf_202_CLK _00693_ VGND VGND VPWR VPWR registers\[5\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_35367_ clknet_leaf_461_CLK _03481_ VGND VGND VPWR VPWR registers\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22332_ registers\[48\]\[47\] registers\[49\]\[47\] registers\[50\]\[47\] registers\[51\]\[47\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__mux4_1
X_25120_ _10817_ registers\[52\]\[41\] _10815_ VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__mux2_1
XFILLER_104_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34318_ clknet_leaf_112_CLK _02432_ VGND VGND VPWR VPWR registers\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35298_ clknet_leaf_473_CLK _03412_ VGND VGND VPWR VPWR registers\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25051_ _10770_ registers\[52\]\[19\] _10752_ VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__mux2_1
X_34249_ clknet_leaf_237_CLK _02363_ VGND VGND VPWR VPWR registers\[33\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_22263_ registers\[52\]\[45\] registers\[53\]\[45\] registers\[54\]\[45\] registers\[55\]\[45\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__mux4_1
XFILLER_247_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24002_ _09542_ registers\[5\]\[13\] _10172_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__mux2_1
X_21214_ _07586_ _07896_ _07897_ _07589_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__a22o_1
XFILLER_145_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22194_ registers\[48\]\[43\] registers\[49\]\[43\] registers\[50\]\[43\] registers\[51\]\[43\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__mux4_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28810_ _12806_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__clkbuf_1
X_21145_ _07305_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29790_ _13352_ VGND VGND VPWR VPWR _13353_ sky130_fd_sc_hd__buf_4
XFILLER_232_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_14__f_CLK clknet_5_7_0_CLK VGND VGND VPWR VPWR clknet_6_14__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_28741_ _11826_ registers\[26\]\[46\] _12763_ VGND VGND VPWR VPWR _12770_ sky130_fd_sc_hd__mux2_1
XFILLER_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21076_ registers\[12\]\[11\] registers\[13\]\[11\] registers\[14\]\[11\] registers\[15\]\[11\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__mux4_1
X_25953_ _10808_ registers\[46\]\[37\] _11263_ VGND VGND VPWR VPWR _11271_ sky130_fd_sc_hd__mux2_1
XFILLER_219_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20027_ _05122_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__buf_4
X_24904_ _09563_ registers\[53\]\[23\] _10680_ VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__mux2_1
X_28672_ _11757_ registers\[26\]\[13\] _12730_ VGND VGND VPWR VPWR _12734_ sky130_fd_sc_hd__mux2_1
X_25884_ _10739_ registers\[46\]\[4\] _11230_ VGND VGND VPWR VPWR _11235_ sky130_fd_sc_hd__mux2_1
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27623_ registers\[34\]\[28\] _10363_ _12173_ VGND VGND VPWR VPWR _12182_ sky130_fd_sc_hd__mux2_1
X_24835_ _10647_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27554_ _12144_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__clkbuf_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _10611_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__clkbuf_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ registers\[56\]\[37\] registers\[57\]\[37\] registers\[58\]\[37\] registers\[59\]\[37\]
+ _08537_ _08327_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__mux4_1
XFILLER_226_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26505_ _11561_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__clkbuf_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23717_ _09529_ registers\[29\]\[7\] _10017_ VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__mux2_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ registers\[12\]\[7\] registers\[13\]\[7\] registers\[14\]\[7\] registers\[15\]\[7\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__mux4_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27485_ _12108_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_215_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24697_ _09628_ registers\[55\]\[54\] _10569_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__mux2_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29224_ _13051_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26436_ _11513_ VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__buf_4
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23648_ _09942_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__buf_4
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29155_ registers\[23\]\[33\] _13004_ _12998_ VGND VGND VPWR VPWR _13005_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_195_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_195_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26367_ _10817_ registers\[43\]\[41\] _11487_ VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__mux2_1
X_23579_ registers\[61\]\[7\] _09672_ _09943_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__mux2_1
XFILLER_126_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16120_ registers\[8\]\[1\] registers\[9\]\[1\] registers\[10\]\[1\] registers\[11\]\[1\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _14633_ sky130_fd_sc_hd__mux4_1
X_28106_ _12436_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25318_ _10858_ registers\[51\]\[61\] _10864_ VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__mux2_1
XFILLER_183_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29086_ net3 VGND VGND VPWR VPWR _12958_ sky130_fd_sc_hd__clkbuf_4
X_26298_ _11452_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16051_ _14564_ VGND VGND VPWR VPWR _14565_ sky130_fd_sc_hd__clkbuf_4
X_28037_ _11797_ registers\[31\]\[32\] _12397_ VGND VGND VPWR VPWR _12400_ sky130_fd_sc_hd__mux2_1
X_25249_ _10789_ registers\[51\]\[28\] _10887_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19810_ _05093_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29988_ _13423_ VGND VGND VPWR VPWR _13457_ sky130_fd_sc_hd__buf_4
XFILLER_81_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16953_ registers\[56\]\[25\] registers\[57\]\[25\] registers\[58\]\[25\] registers\[59\]\[25\]
+ _15409_ _15199_ VGND VGND VPWR VPWR _15442_ sky130_fd_sc_hd__mux4_1
X_19741_ registers\[40\]\[39\] registers\[41\]\[39\] registers\[42\]\[39\] registers\[43\]\[39\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28939_ _12874_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31950_ clknet_leaf_492_CLK _00128_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
X_19672_ registers\[44\]\[37\] registers\[45\]\[37\] registers\[46\]\[37\] registers\[47\]\[37\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__mux4_1
X_16884_ registers\[36\]\[23\] registers\[37\]\[23\] registers\[38\]\[23\] registers\[39\]\[23\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15375_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18623_ registers\[52\]\[7\] registers\[53\]\[7\] registers\[54\]\[7\] registers\[55\]\[7\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__mux4_1
X_30901_ registers\[10\]\[14\] _12964_ _13933_ VGND VGND VPWR VPWR _13938_ sky130_fd_sc_hd__mux2_1
XFILLER_237_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31881_ _14453_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33620_ clknet_leaf_119_CLK _01734_ VGND VGND VPWR VPWR registers\[42\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30832_ _13901_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__clkbuf_1
X_18554_ _05051_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__buf_6
XFILLER_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17505_ _14567_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__clkbuf_4
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33551_ clknet_leaf_147_CLK _01665_ VGND VGND VPWR VPWR registers\[43\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_233_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18485_ registers\[52\]\[3\] registers\[53\]\[3\] registers\[54\]\[3\] registers\[55\]\[3\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__mux4_1
X_30763_ _13865_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1008 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_470 _00162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_481 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32502_ clknet_leaf_329_CLK _00616_ VGND VGND VPWR VPWR registers\[60\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17436_ registers\[20\]\[38\] registers\[21\]\[38\] registers\[22\]\[38\] registers\[23\]\[38\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15912_ sky130_fd_sc_hd__mux4_1
XFILLER_61_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_492 _00166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33482_ clknet_leaf_162_CLK _01596_ VGND VGND VPWR VPWR registers\[45\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30694_ registers\[12\]\[44\] _13027_ _13824_ VGND VGND VPWR VPWR _13829_ sky130_fd_sc_hd__mux2_1
XFILLER_220_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35221_ clknet_leaf_89_CLK _03335_ VGND VGND VPWR VPWR registers\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_28 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32433_ clknet_leaf_386_CLK _00547_ VGND VGND VPWR VPWR registers\[29\]\[35\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_186_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_186_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_39 _00045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _15815_ _15824_ _15835_ _15844_ VGND VGND VPWR VPWR _15845_ sky130_fd_sc_hd__or4_4
XFILLER_158_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19106_ _05159_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__clkbuf_4
X_16318_ _14819_ _14824_ _14525_ VGND VGND VPWR VPWR _14825_ sky130_fd_sc_hd__o21ba_1
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35152_ clknet_leaf_114_CLK _03266_ VGND VGND VPWR VPWR registers\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32364_ clknet_leaf_374_CLK _00478_ VGND VGND VPWR VPWR registers\[61\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298_ _15777_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34103_ clknet_leaf_343_CLK _02217_ VGND VGND VPWR VPWR registers\[35\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_31315_ _14155_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__clkbuf_1
X_19037_ _05069_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__buf_4
X_35083_ clknet_leaf_143_CLK _03197_ VGND VGND VPWR VPWR registers\[20\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_16249_ _14528_ _14756_ _14757_ _14537_ VGND VGND VPWR VPWR _14758_ sky130_fd_sc_hd__a22o_1
X_32295_ clknet_leaf_449_CLK _00409_ VGND VGND VPWR VPWR registers\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xoutput102 net102 VGND VGND VPWR VPWR D1[20] sky130_fd_sc_hd__buf_2
X_34034_ clknet_leaf_357_CLK _02148_ VGND VGND VPWR VPWR registers\[36\]\[36\] sky130_fd_sc_hd__dfxtp_1
Xoutput113 net113 VGND VGND VPWR VPWR D1[30] sky130_fd_sc_hd__buf_2
X_31246_ _14063_ VGND VGND VPWR VPWR _14119_ sky130_fd_sc_hd__buf_4
Xoutput124 net124 VGND VGND VPWR VPWR D1[40] sky130_fd_sc_hd__buf_2
XFILLER_86_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput135 net135 VGND VGND VPWR VPWR D1[50] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR D1[60] sky130_fd_sc_hd__buf_2
Xoutput157 net157 VGND VGND VPWR VPWR D2[12] sky130_fd_sc_hd__buf_2
XFILLER_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput168 net168 VGND VGND VPWR VPWR D2[22] sky130_fd_sc_hd__buf_2
XFILLER_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput179 net179 VGND VGND VPWR VPWR D2[32] sky130_fd_sc_hd__buf_2
XFILLER_130_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31177_ registers\[8\]\[17\] net9 _14075_ VGND VGND VPWR VPWR _14083_ sky130_fd_sc_hd__mux2_1
XFILLER_86_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30128_ registers\[16\]\[32\] _13002_ _13528_ VGND VGND VPWR VPWR _13531_ sky130_fd_sc_hd__mux2_1
X_19939_ _06379_ _06656_ _06657_ _06382_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__a22o_1
XFILLER_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35985_ clknet_leaf_179_CLK _04099_ VGND VGND VPWR VPWR registers\[63\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30059_ _12933_ _11084_ VGND VGND VPWR VPWR _13494_ sky130_fd_sc_hd__nor2_8
Xclkbuf_leaf_110_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_110_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34936_ clknet_leaf_309_CLK _03050_ VGND VGND VPWR VPWR registers\[22\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_22950_ _09562_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21901_ _08462_ _08563_ _08564_ _08467_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__a22o_1
XFILLER_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_8_0_CLK clknet_2_1_0_CLK VGND VGND VPWR VPWR clknet_5_8_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22881_ _09510_ registers\[62\]\[0\] _09515_ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__mux2_1
XFILLER_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34867_ clknet_leaf_412_CLK _02981_ VGND VGND VPWR VPWR registers\[23\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_848 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24620_ _10533_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
X_21832_ _08498_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__buf_6
X_33818_ clknet_leaf_11_CLK _01932_ VGND VGND VPWR VPWR registers\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34798_ clknet_leaf_385_CLK _02912_ VGND VGND VPWR VPWR registers\[24\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24551_ _09619_ registers\[56\]\[50\] _10495_ VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__mux2_1
X_21763_ _08398_ _08407_ _08417_ _08431_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__or4_1
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33749_ clknet_leaf_125_CLK _01863_ VGND VGND VPWR VPWR registers\[40\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20714_ registers\[48\]\[1\] registers\[49\]\[1\] registers\[50\]\[1\] registers\[51\]\[1\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__mux4_1
X_23502_ _09909_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__clkbuf_1
X_27270_ _11995_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_212_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21694_ registers\[36\]\[29\] registers\[37\]\[29\] registers\[38\]\[29\] registers\[39\]\[29\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__mux4_1
X_24482_ _10459_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26221_ _10806_ registers\[44\]\[36\] _11405_ VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__mux2_1
X_20645_ _07287_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__buf_8
X_23433_ _09873_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__clkbuf_1
X_35419_ clknet_leaf_477_CLK _03533_ VGND VGND VPWR VPWR registers\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_177_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_177_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26152_ _10737_ registers\[44\]\[3\] _11372_ VGND VGND VPWR VPWR _11376_ sky130_fd_sc_hd__mux2_1
XFILLER_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23364_ _09835_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
X_20576_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__buf_12
XFILLER_20_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25103_ net30 VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__buf_2
X_22315_ _08761_ _08964_ _08967_ _08764_ VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__a22o_1
XFILLER_109_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23295_ registers\[9\]\[47\] _09791_ _09776_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__mux2_1
XFILLER_152_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26083_ _11339_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29911_ _13416_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22246_ registers\[28\]\[44\] registers\[29\]\[44\] registers\[30\]\[44\] registers\[31\]\[44\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__mux4_1
X_25034_ _10759_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29842_ _13380_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__clkbuf_1
X_22177_ _08761_ _08832_ _08833_ _08764_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__a22o_1
XFILLER_121_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21128_ registers\[32\]\[13\] registers\[33\]\[13\] registers\[34\]\[13\] registers\[35\]\[13\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__mux4_1
X_29773_ registers\[1\]\[56\] _13052_ _13337_ VGND VGND VPWR VPWR _13344_ sky130_fd_sc_hd__mux2_1
XFILLER_191_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26985_ _11839_ registers\[3\]\[52\] _11835_ VGND VGND VPWR VPWR _11840_ sky130_fd_sc_hd__mux2_1
XFILLER_78_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28724_ _11809_ registers\[26\]\[38\] _12752_ VGND VGND VPWR VPWR _12761_ sky130_fd_sc_hd__mux2_1
XFILLER_87_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_101_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_101_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21059_ registers\[40\]\[11\] registers\[41\]\[11\] registers\[42\]\[11\] registers\[43\]\[11\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__mux4_1
X_25936_ _10791_ registers\[46\]\[29\] _11252_ VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__mux2_1
XFILLER_47_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28655_ _11740_ registers\[26\]\[5\] _12719_ VGND VGND VPWR VPWR _12725_ sky130_fd_sc_hd__mux2_1
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25867_ _11225_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27606_ _12150_ VGND VGND VPWR VPWR _12173_ sky130_fd_sc_hd__buf_4
X_24818_ _10638_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28586_ _12688_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__clkbuf_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25798_ _11189_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27537_ _11839_ registers\[35\]\[52\] _12133_ VGND VGND VPWR VPWR _12136_ sky130_fd_sc_hd__mux2_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24749_ _10602_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ registers\[20\]\[63\] registers\[21\]\[63\] registers\[22\]\[63\] registers\[23\]\[63\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux4_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27468_ _12099_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29207_ _12934_ VGND VGND VPWR VPWR _13040_ sky130_fd_sc_hd__buf_4
X_17221_ _15699_ _15702_ _15631_ VGND VGND VPWR VPWR _15703_ sky130_fd_sc_hd__o21ba_1
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26419_ _11516_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_168_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_168_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27399_ _12063_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29138_ net21 VGND VGND VPWR VPWR _12993_ sky130_fd_sc_hd__clkbuf_4
X_17152_ _14597_ VGND VGND VPWR VPWR _15636_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_844 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput15 DW[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 DW[32] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_155_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 DW[42] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_8
X_16103_ _14616_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_4
Xinput48 DW[52] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_8
XFILLER_171_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput59 DW[62] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_16
X_29069_ _12946_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17083_ registers\[20\]\[28\] registers\[21\]\[28\] registers\[22\]\[28\] registers\[23\]\[28\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15569_ sky130_fd_sc_hd__mux4_1
XFILLER_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31100_ _14042_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__clkbuf_1
X_16034_ _14495_ VGND VGND VPWR VPWR _14548_ sky130_fd_sc_hd__buf_12
XFILLER_170_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32080_ clknet_leaf_491_CLK _00022_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31031_ _14006_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_340_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_340_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_123_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17985_ _04548_ _04756_ _04757_ _04552_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__a22o_1
XFILLER_46_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16936_ _14564_ VGND VGND VPWR VPWR _15426_ sky130_fd_sc_hd__clkbuf_4
X_19724_ registers\[0\]\[38\] registers\[1\]\[38\] registers\[2\]\[38\] registers\[3\]\[38\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__mux4_1
X_32982_ clknet_leaf_65_CLK _01096_ VGND VGND VPWR VPWR registers\[52\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35770_ clknet_leaf_287_CLK _03884_ VGND VGND VPWR VPWR registers\[0\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_6_60__f_CLK clknet_5_30_0_CLK VGND VGND VPWR VPWR clknet_6_60__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_226_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34721_ clknet_leaf_8_CLK _02835_ VGND VGND VPWR VPWR registers\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31933_ _14480_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__clkbuf_1
X_16867_ _15144_ _15357_ _15358_ _15147_ VGND VGND VPWR VPWR _15359_ sky130_fd_sc_hd__a22o_1
X_19655_ _05130_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__buf_4
XFILLER_225_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18606_ _05150_ _05361_ _05362_ _05160_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a22o_1
XFILLER_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19586_ _06036_ _06313_ _06314_ _06039_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__a22o_1
X_34652_ clknet_leaf_4_CLK _02766_ VGND VGND VPWR VPWR registers\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_31864_ _14444_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16798_ registers\[16\]\[20\] registers\[17\]\[20\] registers\[18\]\[20\] registers\[19\]\[20\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15292_ sky130_fd_sc_hd__mux4_1
XFILLER_80_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33603_ clknet_leaf_250_CLK _01717_ VGND VGND VPWR VPWR registers\[43\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_18537_ _05292_ _05295_ _05163_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30815_ _13892_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31795_ registers\[59\]\[54\] net50 _14403_ VGND VGND VPWR VPWR _14408_ sky130_fd_sc_hd__mux2_1
X_34583_ clknet_leaf_93_CLK _02697_ VGND VGND VPWR VPWR registers\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18468_ registers\[28\]\[2\] registers\[29\]\[2\] registers\[30\]\[2\] registers\[31\]\[2\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__mux4_1
X_30746_ _13856_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__clkbuf_1
X_33534_ clknet_leaf_274_CLK _01648_ VGND VGND VPWR VPWR registers\[44\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17419_ registers\[52\]\[38\] registers\[53\]\[38\] registers\[54\]\[38\] registers\[55\]\[38\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _15895_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_159_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_159_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33465_ clknet_leaf_280_CLK _01579_ VGND VGND VPWR VPWR registers\[45\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18399_ net82 net81 VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__or2b_4
X_30677_ registers\[12\]\[36\] _13010_ _13813_ VGND VGND VPWR VPWR _13820_ sky130_fd_sc_hd__mux2_1
XFILLER_165_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35204_ clknet_leaf_219_CLK _03318_ VGND VGND VPWR VPWR registers\[18\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_20430_ _06919_ _07132_ _07133_ _06922_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__a22o_1
X_32416_ clknet_leaf_1_CLK _00530_ VGND VGND VPWR VPWR registers\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36184_ clknet_leaf_92_CLK _00065_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
X_33396_ clknet_leaf_346_CLK _01510_ VGND VGND VPWR VPWR registers\[46\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_20361_ _06873_ _07066_ _07067_ _06878_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__a22o_1
X_35135_ clknet_leaf_300_CLK _03249_ VGND VGND VPWR VPWR registers\[1\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32347_ clknet_leaf_55_CLK _00461_ VGND VGND VPWR VPWR registers\[61\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22100_ _07369_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__buf_2
XFILLER_88_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23080_ net88 VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__buf_6
X_35066_ clknet_leaf_309_CLK _03180_ VGND VGND VPWR VPWR registers\[20\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_20292_ _06722_ _06999_ _07000_ _06725_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__a22o_1
XFILLER_162_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32278_ clknet_leaf_86_CLK _00392_ VGND VGND VPWR VPWR registers\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_22031_ _08686_ _08691_ _08416_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__o21ba_1
X_34017_ clknet_leaf_41_CLK _02131_ VGND VGND VPWR VPWR registers\[36\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31229_ _14110_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_331_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_331_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_216_1226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26770_ _11701_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__clkbuf_1
X_35968_ clknet_leaf_231_CLK _04082_ VGND VGND VPWR VPWR registers\[6\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23982_ _10165_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25721_ registers\[48\]\[56\] _10422_ _11141_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__mux2_1
XFILLER_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34919_ clknet_leaf_456_CLK _03033_ VGND VGND VPWR VPWR registers\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22933_ _09550_ registers\[62\]\[17\] _09536_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__mux2_1
XFILLER_229_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35899_ clknet_leaf_301_CLK _04013_ VGND VGND VPWR VPWR registers\[7\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28440_ _11795_ registers\[28\]\[31\] _12610_ VGND VGND VPWR VPWR _12612_ sky130_fd_sc_hd__mux2_1
X_25652_ registers\[48\]\[23\] _10353_ _11108_ VGND VGND VPWR VPWR _11112_ sky130_fd_sc_hd__mux2_1
X_22864_ _07296_ _09498_ _09499_ _07302_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__a22o_1
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24603_ _10524_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28371_ registers\[2\]\[63\] _10436_ _12505_ VGND VGND VPWR VPWR _12575_ sky130_fd_sc_hd__mux2_1
XFILLER_25_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21815_ registers\[8\]\[32\] registers\[9\]\[32\] registers\[10\]\[32\] registers\[11\]\[32\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__mux4_1
X_25583_ registers\[4\]\[56\] _10422_ _11067_ VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_398_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_398_CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22795_ registers\[60\]\[61\] registers\[61\]\[61\] registers\[62\]\[61\] registers\[63\]\[61\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__mux4_1
XFILLER_19_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1071 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27322_ registers\[36\]\[14\] _10334_ _12018_ VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__mux2_1
XFILLER_224_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24534_ _09603_ registers\[56\]\[42\] _10484_ VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__mux2_1
XFILLER_25_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21746_ _08272_ _08413_ _08414_ _08275_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__a22o_1
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27253_ _11986_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24465_ _10450_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
X_21677_ _08272_ _08344_ _08347_ _08275_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__a22o_1
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26204_ _10789_ registers\[44\]\[28\] _11394_ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__mux2_1
X_23416_ _09862_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20628_ _07326_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__buf_6
XFILLER_32_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27184_ _11950_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__clkbuf_1
X_24396_ _10406_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26135_ _11366_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20559_ registers\[8\]\[63\] registers\[9\]\[63\] registers\[10\]\[63\] registers\[11\]\[63\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__mux4_1
X_23347_ _09826_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26066_ _11330_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
X_23278_ registers\[9\]\[42\] _09780_ _09776_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25017_ _10747_ registers\[52\]\[8\] _10731_ VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__mux2_1
X_22229_ _07326_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__buf_6
XFILLER_156_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_322_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_322_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1605 _14581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1616 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29825_ _13371_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1627 _15845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1638 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1649 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17770_ _14543_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__buf_4
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29756_ registers\[1\]\[48\] _13035_ _13326_ VGND VGND VPWR VPWR _13335_ sky130_fd_sc_hd__mux2_1
X_26968_ net42 VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__buf_4
XFILLER_134_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16721_ _14576_ VGND VGND VPWR VPWR _15217_ sky130_fd_sc_hd__buf_6
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25919_ _11253_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28707_ _12718_ VGND VGND VPWR VPWR _12752_ sky130_fd_sc_hd__buf_4
X_29687_ registers\[1\]\[15\] _12966_ _13293_ VGND VGND VPWR VPWR _13299_ sky130_fd_sc_hd__mux2_1
X_26899_ _11781_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_235_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19440_ _05111_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__buf_6
XFILLER_90_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28638_ _12715_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__clkbuf_1
X_16652_ registers\[24\]\[16\] registers\[25\]\[16\] registers\[26\]\[16\] registers\[27\]\[16\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15150_ sky130_fd_sc_hd__mux4_1
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19371_ registers\[0\]\[28\] registers\[1\]\[28\] registers\[2\]\[28\] registers\[3\]\[28\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_389_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_389_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16583_ _14564_ VGND VGND VPWR VPWR _15083_ sky130_fd_sc_hd__buf_4
X_28569_ _12679_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30600_ _09705_ _11010_ VGND VGND VPWR VPWR _13779_ sky130_fd_sc_hd__nor2_8
X_18322_ registers\[48\]\[0\] registers\[49\]\[0\] registers\[50\]\[0\] registers\[51\]\[0\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31580_ registers\[63\]\[16\] net8 _14288_ VGND VGND VPWR VPWR _14295_ sky130_fd_sc_hd__mux2_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ registers\[48\]\[63\] registers\[49\]\[63\] registers\[50\]\[63\] registers\[51\]\[63\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__mux4_1
XFILLER_124_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30531_ _13743_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17204_ registers\[36\]\[32\] registers\[37\]\[32\] registers\[38\]\[32\] registers\[39\]\[32\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15686_ sky130_fd_sc_hd__mux4_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33250_ clknet_leaf_441_CLK _01364_ VGND VGND VPWR VPWR registers\[48\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_30462_ _13706_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18184_ _04950_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32201_ clknet_leaf_375_CLK _00315_ VGND VGND VPWR VPWR registers\[9\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17135_ _15549_ _15617_ _15618_ _15553_ VGND VGND VPWR VPWR _15619_ sky130_fd_sc_hd__a22o_1
XFILLER_129_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33181_ clknet_leaf_474_CLK _01295_ VGND VGND VPWR VPWR registers\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_30393_ _13670_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32132_ clknet_leaf_460_CLK _00049_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfxtp_1
X_17066_ registers\[52\]\[28\] registers\[53\]\[28\] registers\[54\]\[28\] registers\[55\]\[28\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15552_ sky130_fd_sc_hd__mux4_1
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16017_ _14495_ VGND VGND VPWR VPWR _14531_ sky130_fd_sc_hd__buf_12
XFILLER_98_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32063_ clknet_leaf_293_CLK _00241_ VGND VGND VPWR VPWR registers\[62\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_313_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_313_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31014_ _13997_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__clkbuf_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35822_ clknet_leaf_376_CLK _03936_ VGND VGND VPWR VPWR registers\[8\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17968_ _04738_ _04741_ _04644_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__o21ba_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19707_ _06428_ _06431_ _06161_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__o21ba_1
X_35753_ clknet_leaf_458_CLK _03867_ VGND VGND VPWR VPWR registers\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_16919_ _14529_ VGND VGND VPWR VPWR _15409_ sky130_fd_sc_hd__buf_6
X_32965_ clknet_leaf_294_CLK _01079_ VGND VGND VPWR VPWR registers\[53\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17899_ _04653_ _04660_ _04667_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__or4_4
X_34704_ clknet_leaf_118_CLK _02818_ VGND VGND VPWR VPWR registers\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_31916_ _14471_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__clkbuf_1
X_19638_ registers\[56\]\[36\] registers\[57\]\[36\] registers\[58\]\[36\] registers\[59\]\[36\]
+ _06301_ _06091_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__mux4_1
X_35684_ clknet_leaf_465_CLK _03798_ VGND VGND VPWR VPWR registers\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32896_ clknet_leaf_294_CLK _01010_ VGND VGND VPWR VPWR registers\[54\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34635_ clknet_leaf_152_CLK _02749_ VGND VGND VPWR VPWR registers\[27\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31847_ _14435_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19569_ registers\[36\]\[34\] registers\[37\]\[34\] registers\[38\]\[34\] registers\[39\]\[34\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__mux4_1
XFILLER_206_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21600_ registers\[12\]\[26\] registers\[13\]\[26\] registers\[14\]\[26\] registers\[15\]\[26\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__mux4_1
X_22580_ registers\[48\]\[54\] registers\[49\]\[54\] registers\[50\]\[54\] registers\[51\]\[54\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__mux4_1
X_34566_ clknet_leaf_220_CLK _02680_ VGND VGND VPWR VPWR registers\[28\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31778_ registers\[59\]\[46\] net41 _14392_ VGND VGND VPWR VPWR _14399_ sky130_fd_sc_hd__mux2_1
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21531_ registers\[12\]\[24\] registers\[13\]\[24\] registers\[14\]\[24\] registers\[15\]\[24\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__mux4_1
X_33517_ clknet_leaf_345_CLK _01631_ VGND VGND VPWR VPWR registers\[44\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_30729_ registers\[12\]\[61\] _13062_ _13779_ VGND VGND VPWR VPWR _13847_ sky130_fd_sc_hd__mux2_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34497_ clknet_leaf_240_CLK _02611_ VGND VGND VPWR VPWR registers\[2\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36236_ clknet_leaf_122_CLK _00122_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dfxtp_1
X_24250_ registers\[57\]\[1\] _10307_ _10305_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__mux2_1
X_21462_ registers\[8\]\[22\] registers\[9\]\[22\] registers\[10\]\[22\] registers\[11\]\[22\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__mux4_1
X_33448_ clknet_leaf_59_CLK _01562_ VGND VGND VPWR VPWR registers\[45\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20413_ registers\[4\]\[58\] registers\[5\]\[58\] registers\[6\]\[58\] registers\[7\]\[58\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__mux4_1
X_23201_ _09731_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36167_ clknet_leaf_263_CLK _04281_ VGND VGND VPWR VPWR registers\[49\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33379_ clknet_leaf_57_CLK _01493_ VGND VGND VPWR VPWR registers\[46\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_21393_ _07929_ _08070_ _08071_ _07932_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__a22o_1
X_24181_ _10270_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20344_ _06776_ _07049_ _07050_ _06782_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__a22o_1
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35118_ clknet_leaf_389_CLK _03232_ VGND VGND VPWR VPWR registers\[1\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_23132_ _09688_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_36098_ clknet_leaf_266_CLK _04212_ VGND VGND VPWR VPWR registers\[59\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_27940_ registers\[32\]\[50\] _10409_ _12348_ VGND VGND VPWR VPWR _12349_ sky130_fd_sc_hd__mux2_1
X_23063_ _09638_ registers\[62\]\[59\] _09620_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__mux2_1
X_20275_ registers\[36\]\[54\] registers\[37\]\[54\] registers\[38\]\[54\] registers\[39\]\[54\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_304_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_304_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35049_ clknet_leaf_405_CLK _03163_ VGND VGND VPWR VPWR registers\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22014_ _07285_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__clkbuf_4
XTAP_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27871_ _12312_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26822_ _09868_ _10159_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__nand2_8
XTAP_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29610_ _13258_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29541_ _13210_ VGND VGND VPWR VPWR _13222_ sky130_fd_sc_hd__buf_4
XFILLER_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26753_ registers\[40\]\[31\] _10370_ _11691_ VGND VGND VPWR VPWR _11693_ sky130_fd_sc_hd__mux2_1
X_23965_ _10155_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_1
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25704_ registers\[48\]\[48\] _10405_ _11130_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__mux2_1
X_29472_ _09778_ registers\[21\]\[41\] _13184_ VGND VGND VPWR VPWR _13186_ sky130_fd_sc_hd__mux2_1
X_22916_ _09539_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_807 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26684_ _11655_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__clkbuf_1
X_23896_ _10119_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28423_ _11778_ registers\[28\]\[23\] _12599_ VGND VGND VPWR VPWR _12603_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25635_ registers\[48\]\[15\] _10336_ _11097_ VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__mux2_1
X_22847_ _07313_ _09481_ _09482_ _07322_ VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__a22o_1
XFILLER_182_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28354_ _12566_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__clkbuf_1
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25566_ registers\[4\]\[48\] _10405_ _11056_ VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__mux2_1
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22778_ _07343_ _09415_ _09416_ _07353_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__a22o_1
XFILLER_213_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27305_ registers\[36\]\[6\] _10317_ _12007_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__mux2_1
XFILLER_160_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24517_ _09586_ registers\[56\]\[34\] _10473_ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28285_ _12530_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__clkbuf_1
X_21729_ _08391_ _08396_ _08397_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__o21ba_1
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25497_ registers\[4\]\[15\] _10336_ _11023_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__mux2_1
XFILLER_184_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27236_ _11977_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__clkbuf_1
X_24448_ _09517_ registers\[56\]\[1\] _10440_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__mux2_1
XFILLER_184_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27167_ _11941_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24379_ net38 VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_193_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26118_ _10838_ registers\[45\]\[51\] _11356_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__mux2_1
XFILLER_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27098_ _11805_ registers\[38\]\[36\] _11898_ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26049_ _11321_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
X_18940_ _05681_ _05686_ _05483_ _05484_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o211a_2
XFILLER_45_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1402 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1413 _00181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1424 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18871_ registers\[60\]\[14\] registers\[61\]\[14\] registers\[62\]\[14\] registers\[63\]\[14\]
+ _05619_ _05413_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__mux4_1
XTAP_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1435 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1446 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17822_ _04294_ _04598_ _04599_ _04299_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a22o_1
X_29808_ _13362_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1457 _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1468 _05162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1479 _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29739_ _13281_ VGND VGND VPWR VPWR _13326_ sky130_fd_sc_hd__buf_4
X_17753_ _04532_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_4
XTAP_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16704_ registers\[56\]\[18\] registers\[57\]\[18\] registers\[58\]\[18\] registers\[59\]\[18\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15200_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17684_ registers\[40\]\[46\] registers\[41\]\[46\] registers\[42\]\[46\] registers\[43\]\[46\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__mux4_1
X_32750_ clknet_leaf_371_CLK _00864_ VGND VGND VPWR VPWR registers\[56\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31701_ _14358_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__clkbuf_1
X_19423_ _05095_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__buf_4
X_16635_ registers\[60\]\[16\] registers\[61\]\[16\] registers\[62\]\[16\] registers\[63\]\[16\]
+ _15070_ _14864_ VGND VGND VPWR VPWR _15133_ sky130_fd_sc_hd__mux4_1
X_32681_ clknet_leaf_424_CLK _00795_ VGND VGND VPWR VPWR registers\[57\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_34420_ clknet_leaf_416_CLK _02534_ VGND VGND VPWR VPWR registers\[30\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_31632_ _14322_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__clkbuf_1
X_16566_ _14529_ VGND VGND VPWR VPWR _15066_ sky130_fd_sc_hd__buf_6
X_19354_ _06085_ _06088_ _05818_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__o21ba_1
XFILLER_204_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18305_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__clkbuf_8
X_31563_ registers\[63\]\[8\] net63 _14277_ VGND VGND VPWR VPWR _14286_ sky130_fd_sc_hd__mux2_1
X_34351_ clknet_leaf_411_CLK _02465_ VGND VGND VPWR VPWR registers\[31\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_19285_ registers\[56\]\[26\] registers\[57\]\[26\] registers\[58\]\[26\] registers\[59\]\[26\]
+ _05958_ _05748_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__mux4_1
XFILLER_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16497_ registers\[44\]\[12\] registers\[45\]\[12\] registers\[46\]\[12\] registers\[47\]\[12\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _14999_ sky130_fd_sc_hd__mux4_1
X_18236_ registers\[24\]\[62\] registers\[25\]\[62\] registers\[26\]\[62\] registers\[27\]\[62\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__mux4_1
X_33302_ clknet_leaf_122_CLK _01416_ VGND VGND VPWR VPWR registers\[47\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_30514_ _13734_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34282_ clknet_leaf_427_CLK _02396_ VGND VGND VPWR VPWR registers\[32\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31494_ _14249_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33233_ clknet_leaf_74_CLK _01347_ VGND VGND VPWR VPWR registers\[48\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36021_ clknet_leaf_353_CLK _04135_ VGND VGND VPWR VPWR registers\[63\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_30445_ _09806_ registers\[14\]\[54\] _13693_ VGND VGND VPWR VPWR _13698_ sky130_fd_sc_hd__mux2_1
XFILLER_198_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18167_ _14600_ _04932_ _04933_ _14610_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_90_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_90_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17118_ _15581_ _15588_ _15595_ _15602_ VGND VGND VPWR VPWR _15603_ sky130_fd_sc_hd__or4_4
X_33164_ clknet_leaf_168_CLK _01278_ VGND VGND VPWR VPWR registers\[50\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_1045 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18098_ registers\[44\]\[58\] registers\[45\]\[58\] registers\[46\]\[58\] registers\[47\]\[58\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__mux4_1
XFILLER_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30376_ _09702_ registers\[14\]\[21\] _13660_ VGND VGND VPWR VPWR _13662_ sky130_fd_sc_hd__mux2_1
XFILLER_132_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32115_ clknet_leaf_467_CLK _00030_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dfxtp_1
X_17049_ registers\[32\]\[28\] registers\[33\]\[28\] registers\[34\]\[28\] registers\[35\]\[28\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15535_ sky130_fd_sc_hd__mux4_1
X_33095_ clknet_leaf_260_CLK _01209_ VGND VGND VPWR VPWR registers\[51\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_217_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20060_ _06771_ _06774_ _06504_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__o21ba_1
X_32046_ clknet_leaf_370_CLK _00224_ VGND VGND VPWR VPWR registers\[62\]\[32\] sky130_fd_sc_hd__dfxtp_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35805_ clknet_leaf_484_CLK _03919_ VGND VGND VPWR VPWR registers\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33997_ clknet_leaf_172_CLK _02111_ VGND VGND VPWR VPWR registers\[37\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23750_ _10042_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
X_35736_ clknet_leaf_11_CLK _03850_ VGND VGND VPWR VPWR registers\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _07648_ _07650_ _07651_ _07652_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__a22o_1
X_32948_ clknet_leaf_351_CLK _01062_ VGND VGND VPWR VPWR registers\[53\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_226_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22701_ _09338_ _09341_ _09083_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__o21ba_2
XFILLER_183_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23681_ _10004_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__clkbuf_1
X_35667_ clknet_leaf_79_CLK _03781_ VGND VGND VPWR VPWR registers\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _07295_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__buf_4
X_32879_ clknet_leaf_368_CLK _00993_ VGND VGND VPWR VPWR registers\[54\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25420_ _10986_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
X_22632_ _09272_ _09275_ _09116_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34618_ clknet_leaf_184_CLK _02732_ VGND VGND VPWR VPWR registers\[27\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1060 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35598_ clknet_leaf_109_CLK _03712_ VGND VGND VPWR VPWR registers\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25351_ _10950_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__clkbuf_1
X_22563_ registers\[16\]\[53\] registers\[17\]\[53\] registers\[18\]\[53\] registers\[19\]\[53\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34549_ clknet_leaf_414_CLK _02663_ VGND VGND VPWR VPWR registers\[28\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24302_ registers\[57\]\[18\] _10342_ _10326_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__mux2_1
XFILLER_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28070_ _11830_ registers\[31\]\[48\] _12408_ VGND VGND VPWR VPWR _12417_ sky130_fd_sc_hd__mux2_1
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21514_ _08119_ _08187_ _08188_ _08124_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__a22o_1
XFILLER_210_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25282_ _10913_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__clkbuf_1
X_22494_ _09104_ _09140_ _09141_ _09107_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__a22o_1
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27021_ _11863_ _10585_ VGND VGND VPWR VPWR _11864_ sky130_fd_sc_hd__nand2_8
XFILLER_210_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36219_ clknet_leaf_116_CLK _00103_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dfxtp_1
X_24233_ _10297_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21445_ registers\[40\]\[22\] registers\[41\]\[22\] registers\[42\]\[22\] registers\[43\]\[22\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__mux4_1
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_81_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24164_ _10261_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
X_21376_ _08048_ _08053_ _08054_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20327_ registers\[16\]\[55\] registers\[17\]\[55\] registers\[18\]\[55\] registers\[19\]\[55\]
+ _06729_ _06730_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__mux4_1
X_23115_ registers\[39\]\[9\] _09676_ _09658_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__mux2_1
X_24095_ _10224_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28972_ _12891_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20258_ registers\[12\]\[53\] registers\[13\]\[53\] registers\[14\]\[53\] registers\[15\]\[53\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__mux4_1
X_23046_ _09627_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
X_27923_ registers\[32\]\[42\] _10393_ _12337_ VGND VGND VPWR VPWR _12340_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27854_ _12303_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__clkbuf_1
X_20189_ registers\[4\]\[51\] registers\[5\]\[51\] registers\[6\]\[51\] registers\[7\]\[51\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__mux4_1
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26805_ registers\[40\]\[56\] _10422_ _11713_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__mux2_1
XFILLER_218_910 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27785_ _12267_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__clkbuf_1
X_24997_ _10734_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29524_ _13213_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__clkbuf_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26736_ registers\[40\]\[23\] _10353_ _11680_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__mux2_1
X_23948_ _09624_ registers\[60\]\[52\] _10144_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__mux2_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_800 _08936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_811 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_822 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29455_ _09760_ registers\[21\]\[33\] _13173_ VGND VGND VPWR VPWR _13177_ sky130_fd_sc_hd__mux2_1
X_26667_ _10846_ registers\[41\]\[55\] _11641_ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__mux2_1
XANTENNA_833 _09148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23879_ _10110_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_844 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_855 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_205_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16420_ registers\[36\]\[10\] registers\[37\]\[10\] registers\[38\]\[10\] registers\[39\]\[10\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _14924_ sky130_fd_sc_hd__mux4_1
XANTENNA_866 _09335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25618_ registers\[48\]\[7\] _10319_ _11086_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__mux2_1
X_28406_ _11761_ registers\[28\]\[15\] _12588_ VGND VGND VPWR VPWR _12594_ sky130_fd_sc_hd__mux2_1
XFILLER_232_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29386_ _09648_ registers\[21\]\[0\] _13140_ VGND VGND VPWR VPWR _13141_ sky130_fd_sc_hd__mux2_1
XANTENNA_877 _09529_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26598_ _10777_ registers\[41\]\[22\] _11608_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__mux2_1
XANTENNA_888 _09613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_899 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28337_ _12557_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__clkbuf_1
X_16351_ registers\[56\]\[8\] registers\[57\]\[8\] registers\[58\]\[8\] registers\[59\]\[8\]
+ _14723_ _14856_ VGND VGND VPWR VPWR _14857_ sky130_fd_sc_hd__mux4_1
XFILLER_38_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25549_ _11011_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__buf_4
XFILLER_9_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19070_ _05095_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__buf_4
XFILLER_199_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16282_ registers\[60\]\[6\] registers\[61\]\[6\] registers\[62\]\[6\] registers\[63\]\[6\]
+ _14727_ _14544_ VGND VGND VPWR VPWR _14790_ sky130_fd_sc_hd__mux4_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28268_ _12521_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18021_ _04481_ _04791_ _04792_ _04484_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__a22o_1
XFILLER_240_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27219_ _11968_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28199_ _11824_ registers\[30\]\[45\] _12479_ VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_72_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30230_ _13584_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1_0_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_1_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_158_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30161_ registers\[16\]\[48\] _13035_ _13539_ VGND VGND VPWR VPWR _13548_ sky130_fd_sc_hd__mux2_1
XFILLER_126_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19972_ registers\[4\]\[45\] registers\[5\]\[45\] registers\[6\]\[45\] registers\[7\]\[45\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__mux4_1
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18923_ _05647_ _05654_ _05663_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__or4_2
X_30092_ registers\[16\]\[15\] _12966_ _13506_ VGND VGND VPWR VPWR _13512_ sky130_fd_sc_hd__mux2_1
XFILLER_84_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1210 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1221 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1232 _00034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33920_ clknet_leaf_260_CLK _02034_ VGND VGND VPWR VPWR registers\[38\]\[50\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1243 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18854_ registers\[20\]\[13\] registers\[21\]\[13\] registers\[22\]\[13\] registers\[23\]\[13\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__mux4_1
XFILLER_228_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1254 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1265 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1276 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1287 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17805_ _04540_ _04581_ _04582_ _04546_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__a22o_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1298 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33851_ clknet_leaf_301_CLK _01965_ VGND VGND VPWR VPWR registers\[3\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_15997_ _14510_ VGND VGND VPWR VPWR _14511_ sky130_fd_sc_hd__buf_4
X_18785_ _05501_ _05535_ _05536_ _05506_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__a22o_1
XFILLER_83_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32802_ clknet_leaf_443_CLK _00916_ VGND VGND VPWR VPWR registers\[55\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17736_ _15892_ _04514_ _04515_ _15896_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a22o_1
XFILLER_94_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30994_ _13986_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33782_ clknet_leaf_341_CLK _01896_ VGND VGND VPWR VPWR registers\[40\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_35521_ clknet_leaf_236_CLK _03635_ VGND VGND VPWR VPWR registers\[13\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32733_ clknet_leaf_51_CLK _00847_ VGND VGND VPWR VPWR registers\[56\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17667_ _14504_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__buf_4
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19406_ _06031_ _06138_ _06139_ _06034_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__a22o_1
XFILLER_165_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35452_ clknet_leaf_306_CLK _03566_ VGND VGND VPWR VPWR registers\[14\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_16618_ _14947_ _15115_ _15116_ _14950_ VGND VGND VPWR VPWR _15117_ sky130_fd_sc_hd__a22o_1
XFILLER_51_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32664_ clknet_leaf_68_CLK _00778_ VGND VGND VPWR VPWR registers\[57\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_17598_ _15892_ _04380_ _04381_ _15896_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__a22o_1
XFILLER_35_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34403_ clknet_leaf_473_CLK _02517_ VGND VGND VPWR VPWR registers\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19337_ _06036_ _06071_ _06072_ _06039_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__a22o_1
X_31615_ _14313_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__clkbuf_1
X_16549_ _15044_ _15049_ _14945_ VGND VGND VPWR VPWR _15050_ sky130_fd_sc_hd__o21ba_1
XFILLER_147_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35383_ clknet_leaf_320_CLK _03497_ VGND VGND VPWR VPWR registers\[15\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_32595_ clknet_leaf_73_CLK _00709_ VGND VGND VPWR VPWR registers\[58\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34334_ clknet_leaf_492_CLK _02448_ VGND VGND VPWR VPWR registers\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31546_ _14276_ VGND VGND VPWR VPWR _14277_ sky130_fd_sc_hd__buf_4
X_19268_ _06002_ _06005_ _05837_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__o21ba_1
XFILLER_104_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18219_ registers\[36\]\[62\] registers\[37\]\[62\] registers\[38\]\[62\] registers\[39\]\[62\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux4_1
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34265_ clknet_leaf_90_CLK _02379_ VGND VGND VPWR VPWR registers\[32\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_31477_ _09756_ registers\[6\]\[31\] _14239_ VGND VGND VPWR VPWR _14241_ sky130_fd_sc_hd__mux2_1
X_19199_ registers\[12\]\[23\] registers\[13\]\[23\] registers\[14\]\[23\] registers\[15\]\[23\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__mux4_1
XFILLER_157_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_63_CLK sky130_fd_sc_hd__clkbuf_16
X_36004_ clknet_leaf_446_CLK _04118_ VGND VGND VPWR VPWR registers\[63\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_21230_ _07783_ _07911_ _07912_ _07786_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__a22o_1
X_33216_ clknet_leaf_234_CLK _01330_ VGND VGND VPWR VPWR registers\[4\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30428_ _09788_ registers\[14\]\[46\] _13682_ VGND VGND VPWR VPWR _13689_ sky130_fd_sc_hd__mux2_1
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34196_ clknet_leaf_121_CLK _02310_ VGND VGND VPWR VPWR registers\[33\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21161_ _07776_ _07844_ _07845_ _07781_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__a22o_1
X_33147_ clknet_leaf_283_CLK _01261_ VGND VGND VPWR VPWR registers\[50\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_30359_ _09685_ registers\[14\]\[13\] _13649_ VGND VGND VPWR VPWR _13653_ sky130_fd_sc_hd__mux2_1
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20112_ _06717_ _06824_ _06825_ _06720_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__a22o_1
X_21092_ registers\[40\]\[12\] registers\[41\]\[12\] registers\[42\]\[12\] registers\[43\]\[12\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__mux4_1
X_33078_ clknet_leaf_334_CLK _01192_ VGND VGND VPWR VPWR registers\[51\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20043_ _06722_ _06757_ _06758_ _06725_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__a22o_1
X_32029_ clknet_leaf_55_CLK _00207_ VGND VGND VPWR VPWR registers\[62\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_24920_ _10692_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _10655_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23802_ _10069_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27570_ _12154_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__clkbuf_1
X_24782_ _10619_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21994_ _08418_ _08654_ _08655_ _08421_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__a22o_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26521_ _10835_ registers\[42\]\[50\] _11569_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__mux2_1
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35719_ clknet_leaf_155_CLK _03833_ VGND VGND VPWR VPWR registers\[10\]\[57\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_118 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23733_ _10033_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ registers\[44\]\[8\] registers\[45\]\[8\] registers\[46\]\[8\] registers\[47\]\[8\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__mux4_1
XANTENNA_129 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29240_ net58 VGND VGND VPWR VPWR _13062_ sky130_fd_sc_hd__buf_2
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26452_ _11533_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23664_ _09995_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__clkbuf_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ registers\[36\]\[6\] registers\[37\]\[6\] registers\[38\]\[6\] registers\[39\]\[6\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__mux4_1
X_25403_ _10977_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__clkbuf_1
X_22615_ registers\[60\]\[55\] registers\[61\]\[55\] registers\[62\]\[55\] registers\[63\]\[55\]
+ _09227_ _09021_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__mux4_1
X_29171_ _13015_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__clkbuf_1
X_26383_ _10833_ registers\[43\]\[49\] _11487_ VGND VGND VPWR VPWR _11497_ sky130_fd_sc_hd__mux2_1
X_23595_ _09959_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28122_ _12444_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_37__f_CLK clknet_5_18_0_CLK VGND VGND VPWR VPWR clknet_6_37__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_25334_ _10941_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22546_ registers\[56\]\[53\] registers\[57\]\[53\] registers\[58\]\[53\] registers\[59\]\[53\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__mux4_1
XFILLER_122_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28053_ _12363_ VGND VGND VPWR VPWR _12408_ sky130_fd_sc_hd__clkbuf_8
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25265_ _10904_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__clkbuf_1
X_22477_ _09121_ _09124_ _09083_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__o21ba_1
XFILLER_167_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_54_CLK sky130_fd_sc_hd__clkbuf_16
X_27004_ _11852_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_1
X_24216_ _09619_ registers\[58\]\[50\] _10288_ VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21428_ _07924_ _08104_ _08105_ _07927_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__a22o_1
X_25196_ _10868_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24147_ _10252_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21359_ registers\[16\]\[19\] registers\[17\]\[19\] registers\[18\]\[19\] registers\[19\]\[19\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__mux4_1
XFILLER_159_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24078_ _10215_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28955_ _12882_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23029_ _09615_ registers\[62\]\[48\] _09599_ VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__mux2_1
X_27906_ registers\[32\]\[34\] _10376_ _12326_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28886_ _12846_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__clkbuf_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27837_ registers\[32\]\[1\] _10307_ _12293_ VGND VGND VPWR VPWR _12295_ sky130_fd_sc_hd__mux2_1
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18570_ _05304_ _05311_ _05320_ _05327_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or4_4
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27768_ _12258_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__clkbuf_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29507_ _09815_ registers\[21\]\[58\] _13195_ VGND VGND VPWR VPWR _13204_ sky130_fd_sc_hd__mux2_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17521_ registers\[44\]\[41\] registers\[45\]\[41\] registers\[46\]\[41\] registers\[47\]\[41\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__mux4_1
XFILLER_229_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26719_ registers\[40\]\[15\] _10336_ _11669_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__mux2_1
XFILLER_233_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27699_ _12221_ VGND VGND VPWR VPWR _12222_ sky130_fd_sc_hd__buf_6
XFILLER_72_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_630 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_641 _05162_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_652 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ _15884_ _15925_ _15926_ _15890_ VGND VGND VPWR VPWR _15927_ sky130_fd_sc_hd__a22o_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29438_ _09742_ registers\[21\]\[25\] _13162_ VGND VGND VPWR VPWR _13168_ sky130_fd_sc_hd__mux2_1
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_663 _05297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_674 _05724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16403_ _14801_ _14906_ _14907_ _14804_ VGND VGND VPWR VPWR _14908_ sky130_fd_sc_hd__a22o_1
XANTENNA_685 _06224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_696 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17383_ _15549_ _15858_ _15859_ _15553_ VGND VGND VPWR VPWR _15860_ sky130_fd_sc_hd__a22o_1
X_29369_ _13131_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31400_ registers\[7\]\[59\] net55 _14190_ VGND VGND VPWR VPWR _14200_ sky130_fd_sc_hd__mux2_1
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16334_ registers\[16\]\[7\] registers\[17\]\[7\] registers\[18\]\[7\] registers\[19\]\[7\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _14841_ sky130_fd_sc_hd__mux4_1
X_19122_ registers\[60\]\[21\] registers\[61\]\[21\] registers\[62\]\[21\] registers\[63\]\[21\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__mux4_1
X_32380_ clknet_leaf_288_CLK _00494_ VGND VGND VPWR VPWR registers\[61\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31331_ registers\[7\]\[26\] net19 _14157_ VGND VGND VPWR VPWR _14164_ sky130_fd_sc_hd__mux2_1
X_19053_ _05688_ _05795_ _05796_ _05691_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a22o_1
X_16265_ _14588_ _14772_ _14773_ _14598_ VGND VGND VPWR VPWR _14774_ sky130_fd_sc_hd__a22o_1
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_45_CLK sky130_fd_sc_hd__clkbuf_16
X_18004_ _04776_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31262_ _14127_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__clkbuf_1
X_34050_ clknet_leaf_260_CLK _02164_ VGND VGND VPWR VPWR registers\[36\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_16196_ _14701_ _14706_ _14585_ VGND VGND VPWR VPWR _14707_ sky130_fd_sc_hd__o21ba_1
XFILLER_236_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30213_ _13575_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33001_ clknet_leaf_423_CLK _01115_ VGND VGND VPWR VPWR registers\[52\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31193_ _14091_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30144_ _13494_ VGND VGND VPWR VPWR _13539_ sky130_fd_sc_hd__buf_4
X_19955_ registers\[44\]\[45\] registers\[45\]\[45\] registers\[46\]\[45\] registers\[47\]\[45\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__mux4_1
XFILLER_49_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18906_ _05650_ _05653_ _05483_ _05484_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o211a_2
XFILLER_68_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34952_ clknet_leaf_210_CLK _03066_ VGND VGND VPWR VPWR registers\[22\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_30075_ registers\[16\]\[7\] _12949_ _13495_ VGND VGND VPWR VPWR _13503_ sky130_fd_sc_hd__mux2_1
X_19886_ registers\[40\]\[43\] registers\[41\]\[43\] registers\[42\]\[43\] registers\[43\]\[43\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__mux4_1
XANTENNA_1040 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1051 _13423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1062 _13992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33903_ clknet_leaf_356_CLK _02017_ VGND VGND VPWR VPWR registers\[38\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_18837_ registers\[60\]\[13\] registers\[61\]\[13\] registers\[62\]\[13\] registers\[63\]\[13\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__mux4_1
XANTENNA_1073 _14418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34883_ clknet_leaf_204_CLK _02997_ VGND VGND VPWR VPWR registers\[23\]\[53\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1084 _14500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1095 _14524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33834_ clknet_leaf_401_CLK _01948_ VGND VGND VPWR VPWR registers\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18768_ _05404_ _05518_ _05519_ _05410_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__a22o_1
XFILLER_243_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17719_ _04496_ _04499_ _04301_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__o21ba_1
XFILLER_58_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33765_ clknet_leaf_57_CLK _01879_ VGND VGND VPWR VPWR registers\[40\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_30977_ registers\[10\]\[50\] _13039_ _13977_ VGND VGND VPWR VPWR _13978_ sky130_fd_sc_hd__mux2_1
X_18699_ registers\[0\]\[9\] registers\[1\]\[9\] registers\[2\]\[9\] registers\[3\]\[9\]
+ _05112_ _05114_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__mux4_1
X_35504_ clknet_leaf_375_CLK _03618_ VGND VGND VPWR VPWR registers\[13\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_20730_ registers\[28\]\[1\] registers\[29\]\[1\] registers\[30\]\[1\] registers\[31\]\[1\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__mux4_1
X_32716_ clknet_leaf_168_CLK _00830_ VGND VGND VPWR VPWR registers\[57\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33696_ clknet_leaf_33_CLK _01810_ VGND VGND VPWR VPWR registers\[41\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35435_ clknet_leaf_397_CLK _03549_ VGND VGND VPWR VPWR registers\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20661_ registers\[12\]\[0\] registers\[13\]\[0\] registers\[14\]\[0\] registers\[15\]\[0\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__mux4_1
X_32647_ clknet_leaf_262_CLK _00761_ VGND VGND VPWR VPWR registers\[58\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22400_ registers\[36\]\[49\] registers\[37\]\[49\] registers\[38\]\[49\] registers\[39\]\[49\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__mux4_1
XFILLER_51_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20592_ registers\[32\]\[0\] registers\[33\]\[0\] registers\[34\]\[0\] registers\[35\]\[0\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__mux4_1
XFILLER_220_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23380_ registers\[39\]\[43\] _09782_ _09840_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35366_ clknet_leaf_461_CLK _03480_ VGND VGND VPWR VPWR registers\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32578_ clknet_leaf_233_CLK _00692_ VGND VGND VPWR VPWR registers\[5\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1069 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34317_ clknet_leaf_170_CLK _02431_ VGND VGND VPWR VPWR registers\[32\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22331_ registers\[56\]\[47\] registers\[57\]\[47\] registers\[58\]\[47\] registers\[59\]\[47\]
+ _08880_ _08670_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__mux4_1
X_31529_ _09810_ registers\[6\]\[56\] _14261_ VGND VGND VPWR VPWR _14268_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_36_CLK sky130_fd_sc_hd__clkbuf_16
X_35297_ clknet_leaf_479_CLK _03411_ VGND VGND VPWR VPWR registers\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_25050_ net11 VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__buf_2
X_34248_ clknet_leaf_245_CLK _02362_ VGND VGND VPWR VPWR registers\[33\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22262_ registers\[60\]\[45\] registers\[61\]\[45\] registers\[62\]\[45\] registers\[63\]\[45\]
+ _08884_ _08678_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__mux4_1
XFILLER_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24001_ _10175_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
X_21213_ registers\[4\]\[15\] registers\[5\]\[15\] registers\[6\]\[15\] registers\[7\]\[15\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__mux4_1
X_22193_ registers\[56\]\[43\] registers\[57\]\[43\] registers\[58\]\[43\] registers\[59\]\[43\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__mux4_1
X_34179_ clknet_leaf_247_CLK _02293_ VGND VGND VPWR VPWR registers\[34\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21144_ _07303_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__buf_4
XFILLER_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28740_ _12769_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__clkbuf_1
X_25952_ _11270_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
X_21075_ _07581_ _07761_ _07762_ _07584_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__a22o_1
XFILLER_232_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20026_ _05120_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__buf_4
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24903_ _10683_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28671_ _12733_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25883_ _11234_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24834_ _09628_ registers\[54\]\[54\] _10642_ VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__mux2_1
XFILLER_115_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27622_ _12181_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27553_ _11855_ registers\[35\]\[60\] _12077_ VGND VGND VPWR VPWR _12144_ sky130_fd_sc_hd__mux2_1
X_24765_ _09559_ registers\[54\]\[21\] _10609_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__mux2_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _08633_ _08638_ _08397_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__o21ba_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26504_ _10819_ registers\[42\]\[42\] _11558_ VGND VGND VPWR VPWR _11561_ sky130_fd_sc_hd__mux2_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23716_ _10024_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20928_ _07581_ _07618_ _07619_ _07584_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__a22o_1
XFILLER_148_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27484_ _11786_ registers\[35\]\[27\] _12100_ VGND VGND VPWR VPWR _12108_ sky130_fd_sc_hd__mux2_1
X_24696_ _10573_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26435_ _11524_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__clkbuf_1
X_29223_ registers\[23\]\[55\] _13050_ _13040_ VGND VGND VPWR VPWR _13051_ sky130_fd_sc_hd__mux2_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23647_ _09986_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20859_ registers\[12\]\[5\] registers\[13\]\[5\] registers\[14\]\[5\] registers\[15\]\[5\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__mux4_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29154_ net27 VGND VGND VPWR VPWR _13004_ sky130_fd_sc_hd__clkbuf_4
X_26366_ _11488_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23578_ _09950_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
X_28105_ _11728_ registers\[30\]\[0\] _12435_ VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__mux2_1
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25317_ _10931_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22529_ registers\[16\]\[52\] registers\[17\]\[52\] registers\[18\]\[52\] registers\[19\]\[52\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__mux4_1
X_29085_ _12957_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__clkbuf_1
X_26297_ _10747_ registers\[43\]\[8\] _11443_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_27_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_27_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16050_ _14531_ VGND VGND VPWR VPWR _14564_ sky130_fd_sc_hd__buf_12
X_28036_ _12399_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25248_ _10895_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25179_ _10857_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29987_ _13456_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19740_ _06464_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28938_ registers\[24\]\[11\] _10328_ _12872_ VGND VGND VPWR VPWR _12874_ sky130_fd_sc_hd__mux2_1
X_16952_ _15437_ _15440_ _15269_ VGND VGND VPWR VPWR _15441_ sky130_fd_sc_hd__o21ba_1
XFILLER_238_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19671_ _06226_ _06395_ _06396_ _06231_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__a22o_1
X_16883_ registers\[44\]\[23\] registers\[45\]\[23\] registers\[46\]\[23\] registers\[47\]\[23\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15374_ sky130_fd_sc_hd__mux4_1
X_28869_ _12837_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__clkbuf_1
X_18622_ registers\[60\]\[7\] registers\[61\]\[7\] registers\[62\]\[7\] registers\[63\]\[7\]
+ _05276_ _05093_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__mux4_1
X_30900_ _13937_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__clkbuf_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31880_ _09753_ registers\[49\]\[30\] _14452_ VGND VGND VPWR VPWR _14453_ sky130_fd_sc_hd__mux2_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _05307_ _05310_ _05103_ _05105_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__o211a_1
X_30831_ _09786_ registers\[11\]\[45\] _13895_ VGND VGND VPWR VPWR _13901_ sky130_fd_sc_hd__mux2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ registers\[16\]\[40\] registers\[17\]\[40\] registers\[18\]\[40\] registers\[19\]\[40\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__mux4_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33550_ clknet_leaf_147_CLK _01664_ VGND VGND VPWR VPWR registers\[43\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18484_ registers\[60\]\[3\] registers\[61\]\[3\] registers\[62\]\[3\] registers\[63\]\[3\]
+ _05091_ _05093_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__mux4_1
X_30762_ _09683_ registers\[11\]\[12\] _13862_ VGND VGND VPWR VPWR _13865_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_460 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_471 _00163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32501_ clknet_leaf_353_CLK _00615_ VGND VGND VPWR VPWR registers\[60\]\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ registers\[28\]\[38\] registers\[29\]\[38\] registers\[30\]\[38\] registers\[31\]\[38\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15911_ sky130_fd_sc_hd__mux4_1
XANTENNA_482 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33481_ clknet_leaf_255_CLK _01595_ VGND VGND VPWR VPWR registers\[45\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_30693_ _13828_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_493 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35220_ clknet_leaf_93_CLK _03334_ VGND VGND VPWR VPWR registers\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32432_ clknet_leaf_388_CLK _00546_ VGND VGND VPWR VPWR registers\[29\]\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_18 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_29 _00032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _15840_ _15843_ _15645_ VGND VGND VPWR VPWR _15844_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_20__f_CLK clknet_5_10_0_CLK VGND VGND VPWR VPWR clknet_6_20__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19105_ registers\[20\]\[20\] registers\[21\]\[20\] registers\[22\]\[20\] registers\[23\]\[20\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__mux4_1
X_16317_ _14655_ _14820_ _14823_ _14658_ VGND VGND VPWR VPWR _14824_ sky130_fd_sc_hd__a22o_1
X_35151_ clknet_leaf_118_CLK _03265_ VGND VGND VPWR VPWR registers\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17297_ _15751_ _15760_ _15767_ _15776_ VGND VGND VPWR VPWR _15777_ sky130_fd_sc_hd__or4_4
X_32363_ clknet_leaf_421_CLK _00477_ VGND VGND VPWR VPWR registers\[61\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_18_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_18_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34102_ clknet_leaf_343_CLK _02216_ VGND VGND VPWR VPWR registers\[35\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_16248_ registers\[48\]\[5\] registers\[49\]\[5\] registers\[50\]\[5\] registers\[51\]\[5\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14757_ sky130_fd_sc_hd__mux4_1
X_31314_ registers\[7\]\[18\] net10 _14146_ VGND VGND VPWR VPWR _14155_ sky130_fd_sc_hd__mux2_1
X_19036_ _05067_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__buf_4
X_35082_ clknet_leaf_143_CLK _03196_ VGND VGND VPWR VPWR registers\[20\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_32294_ clknet_leaf_450_CLK _00408_ VGND VGND VPWR VPWR registers\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31245_ _14118_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__clkbuf_1
Xoutput103 net103 VGND VGND VPWR VPWR D1[21] sky130_fd_sc_hd__buf_2
X_34033_ clknet_leaf_359_CLK _02147_ VGND VGND VPWR VPWR registers\[36\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_16179_ _14655_ _14688_ _14689_ _14658_ VGND VGND VPWR VPWR _14690_ sky130_fd_sc_hd__a22o_1
Xoutput114 net114 VGND VGND VPWR VPWR D1[31] sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR D1[41] sky130_fd_sc_hd__buf_2
Xoutput136 net136 VGND VGND VPWR VPWR D1[51] sky130_fd_sc_hd__buf_2
Xoutput147 net147 VGND VGND VPWR VPWR D1[61] sky130_fd_sc_hd__buf_2
XFILLER_47_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput158 net158 VGND VGND VPWR VPWR D2[13] sky130_fd_sc_hd__buf_2
XFILLER_138_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31176_ _14082_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__clkbuf_1
Xoutput169 net169 VGND VGND VPWR VPWR D2[23] sky130_fd_sc_hd__buf_2
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30127_ _13530_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__clkbuf_1
X_19938_ registers\[4\]\[44\] registers\[5\]\[44\] registers\[6\]\[44\] registers\[7\]\[44\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__mux4_1
XFILLER_130_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35984_ clknet_leaf_177_CLK _04098_ VGND VGND VPWR VPWR registers\[63\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30058_ _13493_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__clkbuf_1
X_34935_ clknet_leaf_308_CLK _03049_ VGND VGND VPWR VPWR registers\[22\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19869_ registers\[0\]\[42\] registers\[1\]\[42\] registers\[2\]\[42\] registers\[3\]\[42\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__mux4_1
XFILLER_233_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21900_ registers\[32\]\[35\] registers\[33\]\[35\] registers\[34\]\[35\] registers\[35\]\[35\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__mux4_1
X_22880_ _09514_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__buf_4
X_34866_ clknet_leaf_386_CLK _02980_ VGND VGND VPWR VPWR registers\[23\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21831_ _08474_ _08481_ _08488_ _08497_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__or4_1
XFILLER_55_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33817_ clknet_leaf_12_CLK _01931_ VGND VGND VPWR VPWR registers\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34797_ clknet_leaf_384_CLK _02911_ VGND VGND VPWR VPWR registers\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24550_ _10439_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__buf_6
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33748_ clknet_leaf_119_CLK _01862_ VGND VGND VPWR VPWR registers\[40\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_21762_ _08422_ _08429_ _08430_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23501_ _09588_ registers\[19\]\[35\] _09903_ VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__mux2_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20713_ registers\[56\]\[1\] registers\[57\]\[1\] registers\[58\]\[1\] registers\[59\]\[1\]
+ _07315_ _07317_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__mux4_1
XFILLER_12_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24481_ _09550_ registers\[56\]\[17\] _10451_ VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__mux2_1
X_33679_ clknet_leaf_147_CLK _01793_ VGND VGND VPWR VPWR registers\[41\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21693_ registers\[44\]\[29\] registers\[45\]\[29\] registers\[46\]\[29\] registers\[47\]\[29\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__mux4_1
XFILLER_180_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26220_ _11411_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
X_23432_ _09519_ registers\[19\]\[2\] _09870_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__mux2_1
X_35418_ clknet_leaf_13_CLK _03532_ VGND VGND VPWR VPWR registers\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_20644_ _07275_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__buf_4
XFILLER_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26151_ _11375_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35349_ clknet_leaf_78_CLK _03463_ VGND VGND VPWR VPWR registers\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_23363_ registers\[39\]\[35\] _09764_ _09829_ VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__mux2_1
X_20575_ net73 net74 VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__nor2b_4
XFILLER_221_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25102_ _10805_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__clkbuf_1
X_22314_ registers\[16\]\[46\] registers\[17\]\[46\] registers\[18\]\[46\] registers\[19\]\[46\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__mux4_1
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26082_ _10802_ registers\[45\]\[34\] _11334_ VGND VGND VPWR VPWR _11339_ sky130_fd_sc_hd__mux2_1
X_23294_ net42 VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_118_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29910_ registers\[18\]\[57\] _13054_ _13408_ VGND VGND VPWR VPWR _13416_ sky130_fd_sc_hd__mux2_1
XFILLER_192_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25033_ _10758_ registers\[52\]\[13\] _10752_ VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__mux2_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22245_ _08761_ _08898_ _08899_ _08764_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__a22o_1
XFILLER_219_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29841_ registers\[18\]\[24\] _12985_ _13375_ VGND VGND VPWR VPWR _13380_ sky130_fd_sc_hd__mux2_1
X_22176_ registers\[16\]\[42\] registers\[17\]\[42\] registers\[18\]\[42\] registers\[19\]\[42\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__mux4_1
XFILLER_105_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21127_ registers\[40\]\[13\] registers\[41\]\[13\] registers\[42\]\[13\] registers\[43\]\[13\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__mux4_1
X_29772_ _13343_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26984_ net48 VGND VGND VPWR VPWR _11839_ sky130_fd_sc_hd__buf_4
XFILLER_232_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_247_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28723_ _12760_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__clkbuf_1
X_21058_ _07746_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
X_25935_ _11261_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20009_ _06722_ _06723_ _06724_ _06725_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__a22o_1
XFILLER_115_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25866_ _10856_ registers\[47\]\[60\] _11158_ VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__mux2_1
X_28654_ _12724_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24817_ _09611_ registers\[54\]\[46\] _10631_ VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__mux2_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27605_ _12172_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25797_ _10787_ registers\[47\]\[27\] _11181_ VGND VGND VPWR VPWR _11189_ sky130_fd_sc_hd__mux2_1
X_28585_ _11805_ registers\[27\]\[36\] _12681_ VGND VGND VPWR VPWR _12688_ sky130_fd_sc_hd__mux2_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27536_ _12135_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__clkbuf_1
X_24748_ _09542_ registers\[54\]\[13\] _10598_ VGND VGND VPWR VPWR _10602_ sky130_fd_sc_hd__mux2_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27467_ _11769_ registers\[35\]\[19\] _12089_ VGND VGND VPWR VPWR _12099_ sky130_fd_sc_hd__mux2_1
X_24679_ _10564_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29206_ net46 VGND VGND VPWR VPWR _13039_ sky130_fd_sc_hd__clkbuf_4
X_17220_ _15487_ _15700_ _15701_ _15490_ VGND VGND VPWR VPWR _15702_ sky130_fd_sc_hd__a22o_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26418_ _10733_ registers\[42\]\[1\] _11514_ VGND VGND VPWR VPWR _11516_ sky130_fd_sc_hd__mux2_1
XFILLER_230_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27398_ registers\[36\]\[50\] _10409_ _12062_ VGND VGND VPWR VPWR _12063_ sky130_fd_sc_hd__mux2_1
XFILLER_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_243_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17151_ registers\[16\]\[30\] registers\[17\]\[30\] registers\[18\]\[30\] registers\[19\]\[30\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15635_ sky130_fd_sc_hd__mux4_1
X_29137_ _12992_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__clkbuf_1
X_26349_ _11479_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 DW[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_4
XFILLER_35_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 DW[33] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
X_16102_ _14526_ _14557_ _14586_ _14615_ VGND VGND VPWR VPWR _14616_ sky130_fd_sc_hd__or4_2
XFILLER_156_856 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput38 DW[43] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
XFILLER_183_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29068_ registers\[23\]\[5\] _12945_ _12935_ VGND VGND VPWR VPWR _12946_ sky130_fd_sc_hd__mux2_1
Xinput49 DW[53] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_8
X_17082_ registers\[28\]\[28\] registers\[29\]\[28\] registers\[30\]\[28\] registers\[31\]\[28\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15568_ sky130_fd_sc_hd__mux4_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16033_ _14546_ VGND VGND VPWR VPWR _14547_ sky130_fd_sc_hd__buf_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28019_ _12390_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31030_ registers\[0\]\[11\] _12958_ _14004_ VGND VGND VPWR VPWR _14006_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17984_ registers\[52\]\[54\] registers\[53\]\[54\] registers\[54\]\[54\] registers\[55\]\[54\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__mux4_1
XFILLER_112_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19723_ registers\[8\]\[38\] registers\[9\]\[38\] registers\[10\]\[38\] registers\[11\]\[38\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux4_1
X_16935_ _14562_ VGND VGND VPWR VPWR _15425_ sky130_fd_sc_hd__buf_6
XFILLER_81_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32981_ clknet_leaf_64_CLK _01095_ VGND VGND VPWR VPWR registers\[52\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34720_ clknet_leaf_9_CLK _02834_ VGND VGND VPWR VPWR registers\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31932_ _09808_ registers\[49\]\[55\] _14474_ VGND VGND VPWR VPWR _14480_ sky130_fd_sc_hd__mux2_1
X_19654_ registers\[4\]\[36\] registers\[5\]\[36\] registers\[6\]\[36\] registers\[7\]\[36\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__mux4_1
X_16866_ registers\[4\]\[22\] registers\[5\]\[22\] registers\[6\]\[22\] registers\[7\]\[22\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15358_ sky130_fd_sc_hd__mux4_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_7_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18605_ registers\[20\]\[6\] registers\[21\]\[6\] registers\[22\]\[6\] registers\[23\]\[6\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__mux4_1
XFILLER_203_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34651_ clknet_leaf_20_CLK _02765_ VGND VGND VPWR VPWR registers\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19585_ registers\[4\]\[34\] registers\[5\]\[34\] registers\[6\]\[34\] registers\[7\]\[34\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__mux4_1
X_31863_ _09717_ registers\[49\]\[22\] _14441_ VGND VGND VPWR VPWR _14444_ sky130_fd_sc_hd__mux2_1
X_16797_ registers\[24\]\[20\] registers\[25\]\[20\] registers\[26\]\[20\] registers\[27\]\[20\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15291_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33602_ clknet_leaf_248_CLK _01716_ VGND VGND VPWR VPWR registers\[43\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_248_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18536_ _05150_ _05293_ _05294_ _05160_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30814_ _09769_ registers\[11\]\[37\] _13884_ VGND VGND VPWR VPWR _13892_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34582_ clknet_leaf_88_CLK _02696_ VGND VGND VPWR VPWR registers\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31794_ _14407_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33533_ clknet_leaf_274_CLK _01647_ VGND VGND VPWR VPWR registers\[44\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30745_ _09666_ registers\[11\]\[4\] _13851_ VGND VGND VPWR VPWR _13856_ sky130_fd_sc_hd__mux2_1
X_18467_ _05152_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__buf_6
XFILLER_221_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_290 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17418_ registers\[60\]\[38\] registers\[61\]\[38\] registers\[62\]\[38\] registers\[63\]\[38\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _15894_ sky130_fd_sc_hd__mux4_1
X_33464_ clknet_leaf_339_CLK _01578_ VGND VGND VPWR VPWR registers\[45\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_18398_ _05150_ _05154_ _05158_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__a22o_1
X_30676_ _13819_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35203_ clknet_leaf_223_CLK _03317_ VGND VGND VPWR VPWR registers\[18\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32415_ clknet_leaf_1_CLK _00529_ VGND VGND VPWR VPWR registers\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_36183_ clknet_leaf_93_CLK _00127_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dfxtp_1
X_17349_ registers\[0\]\[36\] registers\[1\]\[36\] registers\[2\]\[36\] registers\[3\]\[36\]
+ _15624_ _15625_ VGND VGND VPWR VPWR _15827_ sky130_fd_sc_hd__mux4_1
X_33395_ clknet_leaf_346_CLK _01509_ VGND VGND VPWR VPWR registers\[46\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35134_ clknet_leaf_299_CLK _03248_ VGND VGND VPWR VPWR registers\[1\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20360_ registers\[20\]\[56\] registers\[21\]\[56\] registers\[22\]\[56\] registers\[23\]\[56\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__mux4_1
XFILLER_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32346_ clknet_leaf_53_CLK _00460_ VGND VGND VPWR VPWR registers\[61\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19019_ _05688_ _05762_ _05763_ _05691_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__a22o_1
X_20291_ registers\[4\]\[54\] registers\[5\]\[54\] registers\[6\]\[54\] registers\[7\]\[54\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__mux4_1
XFILLER_175_1219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35065_ clknet_leaf_308_CLK _03179_ VGND VGND VPWR VPWR registers\[20\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_32277_ clknet_leaf_89_CLK _00391_ VGND VGND VPWR VPWR registers\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_22030_ _08615_ _08687_ _08690_ _08618_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__a22o_1
X_34016_ clknet_leaf_40_CLK _02130_ VGND VGND VPWR VPWR registers\[36\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_31228_ registers\[8\]\[41\] net36 _14108_ VGND VGND VPWR VPWR _14110_ sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31159_ _14073_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23981_ _09521_ registers\[5\]\[3\] _10161_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__mux2_1
X_35967_ clknet_leaf_200_CLK _04081_ VGND VGND VPWR VPWR registers\[6\]\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25720_ _11147_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22932_ net9 VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__buf_4
X_34918_ clknet_leaf_448_CLK _03032_ VGND VGND VPWR VPWR registers\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35898_ clknet_leaf_302_CLK _04012_ VGND VGND VPWR VPWR registers\[7\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25651_ _11111_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
X_22863_ registers\[4\]\[63\] registers\[5\]\[63\] registers\[6\]\[63\] registers\[7\]\[63\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__mux4_1
X_34849_ clknet_leaf_489_CLK _02963_ VGND VGND VPWR VPWR registers\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_1359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24602_ _09533_ registers\[55\]\[9\] _10514_ VGND VGND VPWR VPWR _10524_ sky130_fd_sc_hd__mux2_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28370_ _12574_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__clkbuf_1
X_21814_ _08477_ _08480_ _08405_ _08406_ VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__o211a_1
X_25582_ _11073_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
X_22794_ _07372_ _09430_ _09431_ _07382_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__a22o_1
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27321_ _12022_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__clkbuf_1
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24533_ _10486_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21745_ registers\[4\]\[30\] registers\[5\]\[30\] registers\[6\]\[30\] registers\[7\]\[30\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__mux4_1
XFILLER_184_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27252_ _11824_ registers\[37\]\[45\] _11980_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__mux2_1
X_24464_ _09533_ registers\[56\]\[9\] _10440_ VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__mux2_1
XFILLER_212_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21676_ registers\[4\]\[28\] registers\[5\]\[28\] registers\[6\]\[28\] registers\[7\]\[28\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__mux4_1
XFILLER_71_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26203_ _11402_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
X_23415_ registers\[39\]\[60\] _09819_ _09657_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__mux2_1
XFILLER_196_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20627_ _07277_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__buf_12
XFILLER_137_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27183_ _11755_ registers\[37\]\[12\] _11947_ VGND VGND VPWR VPWR _11950_ sky130_fd_sc_hd__mux2_1
X_24395_ registers\[57\]\[48\] _10405_ _10389_ VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__mux2_1
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26134_ _10854_ registers\[45\]\[59\] _11356_ VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__mux2_1
XFILLER_165_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23346_ registers\[9\]\[63\] _09825_ _09708_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__mux2_1
XFILLER_164_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20558_ _07254_ _07257_ _05102_ _05104_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__o211a_1
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26065_ _10785_ registers\[45\]\[26\] _11323_ VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__mux2_1
XFILLER_152_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23277_ net37 VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__buf_4
X_20489_ registers\[36\]\[61\] registers\[37\]\[61\] registers\[38\]\[61\] registers\[39\]\[61\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__mux4_1
XFILLER_238_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25016_ net63 VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__buf_4
X_22228_ _08669_ _08881_ _08882_ _08675_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__a22o_1
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1606 _14581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29824_ registers\[18\]\[16\] _12968_ _13364_ VGND VGND VPWR VPWR _13371_ sky130_fd_sc_hd__mux2_1
XANTENNA_1617 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22159_ _08812_ _08813_ _08814_ _08815_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__a22o_1
XANTENNA_1628 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1639 _00026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29755_ _13334_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__clkbuf_1
XTAP_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26967_ _11827_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__clkbuf_1
XTAP_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16720_ registers\[12\]\[18\] registers\[13\]\[18\] registers\[14\]\[18\] registers\[15\]\[18\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15216_ sky130_fd_sc_hd__mux4_1
X_28706_ _12751_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__clkbuf_1
X_25918_ _10772_ registers\[46\]\[20\] _11252_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__mux2_1
XFILLER_235_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29686_ _13298_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__clkbuf_1
X_26898_ _11780_ registers\[3\]\[24\] _11772_ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__mux2_1
X_28637_ _11857_ registers\[27\]\[61\] _12647_ VGND VGND VPWR VPWR _12715_ sky130_fd_sc_hd__mux2_1
X_16651_ _15143_ _15148_ _14945_ VGND VGND VPWR VPWR _15149_ sky130_fd_sc_hd__o21ba_1
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25849_ _11216_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19370_ registers\[8\]\[28\] registers\[9\]\[28\] registers\[10\]\[28\] registers\[11\]\[28\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__mux4_1
X_16582_ _14562_ VGND VGND VPWR VPWR _15082_ sky130_fd_sc_hd__buf_6
X_28568_ _11788_ registers\[27\]\[28\] _12670_ VGND VGND VPWR VPWR _12679_ sky130_fd_sc_hd__mux2_1
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18321_ _05045_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27519_ _12126_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__clkbuf_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28499_ _12642_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18252_ registers\[56\]\[63\] registers\[57\]\[63\] registers\[58\]\[63\] registers\[59\]\[63\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux4_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30530_ _09753_ registers\[13\]\[30\] _13742_ VGND VGND VPWR VPWR _13743_ sky130_fd_sc_hd__mux2_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17203_ registers\[44\]\[32\] registers\[45\]\[32\] registers\[46\]\[32\] registers\[47\]\[32\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15685_ sky130_fd_sc_hd__mux4_1
X_30461_ _09823_ registers\[14\]\[62\] _13637_ VGND VGND VPWR VPWR _13706_ sky130_fd_sc_hd__mux2_1
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18183_ _04928_ _04935_ _04942_ _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__or4_4
XFILLER_50_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32200_ clknet_leaf_376_CLK _00314_ VGND VGND VPWR VPWR registers\[9\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_17134_ registers\[52\]\[30\] registers\[53\]\[30\] registers\[54\]\[30\] registers\[55\]\[30\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15618_ sky130_fd_sc_hd__mux4_1
XFILLER_141_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30392_ _09751_ registers\[14\]\[29\] _13660_ VGND VGND VPWR VPWR _13670_ sky130_fd_sc_hd__mux2_1
X_33180_ clknet_leaf_476_CLK _01294_ VGND VGND VPWR VPWR registers\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_7_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_7_0_CLK sky130_fd_sc_hd__clkbuf_8
X_32131_ clknet_leaf_461_CLK _00048_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfxtp_1
X_17065_ registers\[60\]\[28\] registers\[61\]\[28\] registers\[62\]\[28\] registers\[63\]\[28\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15551_ sky130_fd_sc_hd__mux4_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16016_ _14529_ VGND VGND VPWR VPWR _14530_ sky130_fd_sc_hd__buf_12
XFILLER_100_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32062_ clknet_leaf_292_CLK _00240_ VGND VGND VPWR VPWR registers\[62\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31013_ registers\[0\]\[3\] _12941_ _13993_ VGND VGND VPWR VPWR _13997_ sky130_fd_sc_hd__mux2_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_930 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35821_ clknet_leaf_391_CLK _03935_ VGND VGND VPWR VPWR registers\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17967_ _04637_ _04739_ _04740_ _04642_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__a22o_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_670 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19706_ _06233_ _06429_ _06430_ _06236_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__a22o_1
X_35752_ clknet_leaf_457_CLK _03866_ VGND VGND VPWR VPWR registers\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16918_ _15404_ _15407_ _15269_ VGND VGND VPWR VPWR _15408_ sky130_fd_sc_hd__o21ba_1
X_32964_ clknet_leaf_201_CLK _01078_ VGND VGND VPWR VPWR registers\[53\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_17898_ _04670_ _04673_ _04644_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34703_ clknet_leaf_118_CLK _02817_ VGND VGND VPWR VPWR registers\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31915_ _09791_ registers\[49\]\[47\] _14463_ VGND VGND VPWR VPWR _14471_ sky130_fd_sc_hd__mux2_1
XFILLER_26_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19637_ _06360_ _06363_ _06161_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__o21ba_1
X_35683_ clknet_leaf_466_CLK _03797_ VGND VGND VPWR VPWR registers\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_16849_ _14539_ VGND VGND VPWR VPWR _15341_ sky130_fd_sc_hd__buf_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32895_ clknet_leaf_292_CLK _01009_ VGND VGND VPWR VPWR registers\[54\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34634_ clknet_leaf_152_CLK _02748_ VGND VGND VPWR VPWR registers\[27\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31846_ _09687_ registers\[49\]\[14\] _14430_ VGND VGND VPWR VPWR _14435_ sky130_fd_sc_hd__mux2_1
X_19568_ registers\[44\]\[34\] registers\[45\]\[34\] registers\[46\]\[34\] registers\[47\]\[34\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__mux4_1
XFILLER_59_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18519_ registers\[52\]\[4\] registers\[53\]\[4\] registers\[54\]\[4\] registers\[55\]\[4\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__mux4_1
X_34565_ clknet_leaf_221_CLK _02679_ VGND VGND VPWR VPWR registers\[28\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31777_ _14398_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__clkbuf_1
X_19499_ registers\[32\]\[32\] registers\[33\]\[32\] registers\[34\]\[32\] registers\[35\]\[32\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__mux4_1
XFILLER_94_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_885 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21530_ _07924_ _08203_ _08204_ _07927_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__a22o_1
X_33516_ clknet_leaf_345_CLK _01630_ VGND VGND VPWR VPWR registers\[44\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_30728_ _13846_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__clkbuf_1
X_34496_ clknet_leaf_240_CLK _02610_ VGND VGND VPWR VPWR registers\[2\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36235_ clknet_leaf_121_CLK _00121_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33447_ clknet_leaf_60_CLK _01561_ VGND VGND VPWR VPWR registers\[45\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_21461_ _08134_ _08137_ _08062_ _08063_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__o211a_1
XFILLER_194_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30659_ _13810_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23200_ registers\[39\]\[23\] _09730_ _09700_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__mux2_1
X_20412_ registers\[12\]\[58\] registers\[13\]\[58\] registers\[14\]\[58\] registers\[15\]\[58\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__mux4_1
XFILLER_105_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36166_ clknet_leaf_262_CLK _04280_ VGND VGND VPWR VPWR registers\[49\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24180_ _09584_ registers\[58\]\[33\] _10266_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__mux2_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33378_ clknet_leaf_57_CLK _01492_ VGND VGND VPWR VPWR registers\[46\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_21392_ registers\[4\]\[20\] registers\[5\]\[20\] registers\[6\]\[20\] registers\[7\]\[20\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__mux4_1
XFILLER_147_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35117_ clknet_leaf_388_CLK _03231_ VGND VGND VPWR VPWR registers\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_23131_ registers\[39\]\[14\] _09687_ _09679_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__mux2_1
XFILLER_107_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32329_ clknet_leaf_155_CLK _00443_ VGND VGND VPWR VPWR registers\[19\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_20343_ registers\[48\]\[56\] registers\[49\]\[56\] registers\[50\]\[56\] registers\[51\]\[56\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__mux4_1
X_36097_ clknet_leaf_267_CLK _04211_ VGND VGND VPWR VPWR registers\[59\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_1196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23062_ net55 VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__clkbuf_4
X_35048_ clknet_leaf_457_CLK _03162_ VGND VGND VPWR VPWR registers\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_20274_ registers\[44\]\[54\] registers\[45\]\[54\] registers\[46\]\[54\] registers\[47\]\[54\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__mux4_1
XFILLER_150_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22013_ registers\[48\]\[38\] registers\[49\]\[38\] registers\[50\]\[38\] registers\[51\]\[38\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__mux4_1
XTAP_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27870_ registers\[32\]\[17\] _10340_ _12304_ VGND VGND VPWR VPWR _12312_ sky130_fd_sc_hd__mux2_1
XTAP_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26821_ net1 VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__clkbuf_4
XTAP_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29540_ _13221_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__clkbuf_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23964_ _09640_ registers\[60\]\[60\] _10088_ VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26752_ _11692_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__clkbuf_1
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1085 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25703_ _11138_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
X_22915_ _09538_ registers\[62\]\[11\] _09536_ VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__mux2_1
X_26683_ _10862_ registers\[41\]\[63\] _11585_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__mux2_1
X_29471_ _13185_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23895_ _09571_ registers\[60\]\[27\] _10111_ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__mux2_1
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28422_ _12602_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_1
X_22846_ registers\[32\]\[63\] registers\[33\]\[63\] registers\[34\]\[63\] registers\[35\]\[63\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__mux4_1
X_25634_ _11102_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28353_ registers\[2\]\[54\] _10418_ _12561_ VGND VGND VPWR VPWR _12566_ sky130_fd_sc_hd__mux2_1
X_25565_ _11064_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22777_ registers\[16\]\[60\] registers\[17\]\[60\] registers\[18\]\[60\] registers\[19\]\[60\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__mux4_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_240_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_240_CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27304_ _12013_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__clkbuf_1
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24516_ _10477_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
X_21728_ _07309_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__clkbuf_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28284_ registers\[2\]\[21\] _10349_ _12528_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__mux2_1
X_25496_ _11028_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24447_ _10441_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27235_ _11807_ registers\[37\]\[37\] _11969_ VGND VGND VPWR VPWR _11977_ sky130_fd_sc_hd__mux2_1
X_21659_ _07328_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__clkbuf_8
XFILLER_71_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27166_ _11738_ registers\[37\]\[4\] _11936_ VGND VGND VPWR VPWR _11941_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24378_ _10394_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26117_ _11357_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
X_23329_ _09814_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27097_ _11904_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26048_ _10768_ registers\[45\]\[18\] _11312_ VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__mux2_1
XFILLER_106_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1403 _00173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18870_ _05090_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__buf_6
XTAP_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1414 _00181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1425 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1436 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17821_ registers\[20\]\[49\] registers\[21\]\[49\] registers\[22\]\[49\] registers\[23\]\[49\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__mux4_1
XFILLER_132_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29807_ registers\[18\]\[8\] _12951_ _13353_ VGND VGND VPWR VPWR _13362_ sky130_fd_sc_hd__mux2_1
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1447 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1458 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1469 _05289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27999_ _11759_ registers\[31\]\[14\] _12375_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__mux2_1
XFILLER_58_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17752_ _04510_ _04517_ _04524_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__or4_2
X_29738_ _13325_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__clkbuf_1
XTAP_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ _14531_ VGND VGND VPWR VPWR _15199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_236_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29669_ _13289_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__clkbuf_1
X_17683_ _04464_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_208_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31700_ registers\[59\]\[9\] net64 _14348_ VGND VGND VPWR VPWR _14358_ sky130_fd_sc_hd__mux2_1
X_19422_ _05883_ _06153_ _06154_ _05888_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a22o_1
X_16634_ _14855_ _15130_ _15131_ _14861_ VGND VGND VPWR VPWR _15132_ sky130_fd_sc_hd__a22o_1
X_32680_ clknet_leaf_436_CLK _00794_ VGND VGND VPWR VPWR registers\[57\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19353_ _05890_ _06086_ _06087_ _05893_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__a22o_1
X_31631_ registers\[63\]\[40\] net35 _14321_ VGND VGND VPWR VPWR _14322_ sky130_fd_sc_hd__mux2_1
X_16565_ _15061_ _15064_ _14926_ VGND VGND VPWR VPWR _15065_ sky130_fd_sc_hd__o21ba_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_231_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_231_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18304_ _05041_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__buf_12
X_34350_ clknet_leaf_386_CLK _02464_ VGND VGND VPWR VPWR registers\[31\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_31562_ _14285_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__clkbuf_1
X_19284_ _06017_ _06020_ _05818_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__o21ba_1
X_16496_ _14539_ VGND VGND VPWR VPWR _14998_ sky130_fd_sc_hd__clkbuf_4
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33301_ clknet_leaf_123_CLK _01415_ VGND VGND VPWR VPWR registers\[47\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18235_ _04996_ _04999_ _14584_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o21ba_1
X_30513_ _09717_ registers\[13\]\[22\] _13731_ VGND VGND VPWR VPWR _13734_ sky130_fd_sc_hd__mux2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34281_ clknet_leaf_427_CLK _02395_ VGND VGND VPWR VPWR registers\[32\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31493_ _09773_ registers\[6\]\[39\] _14239_ VGND VGND VPWR VPWR _14249_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36020_ clknet_leaf_324_CLK _04134_ VGND VGND VPWR VPWR registers\[63\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_33232_ clknet_leaf_75_CLK _01346_ VGND VGND VPWR VPWR registers\[48\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_30444_ _13697_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__clkbuf_1
X_18166_ registers\[52\]\[60\] registers\[53\]\[60\] registers\[54\]\[60\] registers\[55\]\[60\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__mux4_1
XFILLER_156_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ _15598_ _15601_ _15302_ VGND VGND VPWR VPWR _15602_ sky130_fd_sc_hd__o21ba_1
XFILLER_102_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33163_ clknet_leaf_164_CLK _01277_ VGND VGND VPWR VPWR registers\[50\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18097_ _04676_ _04864_ _04865_ _04681_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a22o_1
X_30375_ _13661_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32114_ clknet_leaf_467_CLK _00029_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dfxtp_1
X_17048_ registers\[40\]\[28\] registers\[41\]\[28\] registers\[42\]\[28\] registers\[43\]\[28\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15534_ sky130_fd_sc_hd__mux4_1
X_33094_ clknet_leaf_263_CLK _01208_ VGND VGND VPWR VPWR registers\[51\]\[56\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_298_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_298_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32045_ clknet_leaf_374_CLK _00223_ VGND VGND VPWR VPWR registers\[62\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ registers\[36\]\[18\] registers\[37\]\[18\] registers\[38\]\[18\] registers\[39\]\[18\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__mux4_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35804_ clknet_leaf_16_CLK _03918_ VGND VGND VPWR VPWR registers\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_33996_ clknet_leaf_168_CLK _02110_ VGND VGND VPWR VPWR registers\[37\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35735_ clknet_leaf_81_CLK _03849_ VGND VGND VPWR VPWR registers\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20961_ _07301_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32947_ clknet_leaf_355_CLK _01061_ VGND VGND VPWR VPWR registers\[53\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22700_ _09155_ _09339_ _09340_ _09158_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_470_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_470_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23680_ registers\[61\]\[55\] _09808_ _09998_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__mux2_1
X_35666_ clknet_leaf_106_CLK _03780_ VGND VGND VPWR VPWR registers\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20892_ _07581_ _07582_ _07583_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__a22o_1
X_32878_ clknet_leaf_368_CLK _00992_ VGND VGND VPWR VPWR registers\[54\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22631_ _09109_ _09273_ _09274_ _09114_ VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__a22o_1
X_34617_ clknet_leaf_428_CLK _02731_ VGND VGND VPWR VPWR registers\[27\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31829_ _09670_ registers\[49\]\[6\] _14419_ VGND VGND VPWR VPWR _14426_ sky130_fd_sc_hd__mux2_1
X_35597_ clknet_leaf_145_CLK _03711_ VGND VGND VPWR VPWR registers\[12\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_222_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_222_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25350_ _10754_ registers\[50\]\[11\] _10948_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__mux2_1
X_22562_ registers\[24\]\[53\] registers\[25\]\[53\] registers\[26\]\[53\] registers\[27\]\[53\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__mux4_1
XFILLER_210_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34548_ clknet_leaf_415_CLK _02662_ VGND VGND VPWR VPWR registers\[28\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_222_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24301_ net10 VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__buf_4
X_21513_ registers\[32\]\[24\] registers\[33\]\[24\] registers\[34\]\[24\] registers\[35\]\[24\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__mux4_1
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25281_ _10821_ registers\[51\]\[43\] _10909_ VGND VGND VPWR VPWR _10913_ sky130_fd_sc_hd__mux2_1
X_22493_ registers\[16\]\[51\] registers\[17\]\[51\] registers\[18\]\[51\] registers\[19\]\[51\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__mux4_1
X_34479_ clknet_leaf_377_CLK _02593_ VGND VGND VPWR VPWR registers\[2\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_27020_ _09649_ _09650_ _09651_ VGND VGND VPWR VPWR _11863_ sky130_fd_sc_hd__nor3b_4
X_36218_ clknet_leaf_116_CLK _00102_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dfxtp_1
X_24232_ _09636_ registers\[58\]\[58\] _10288_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__mux2_1
XFILLER_33_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21444_ _07281_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__buf_4
XFILLER_147_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24163_ _09567_ registers\[58\]\[25\] _10255_ VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__mux2_1
X_36149_ clknet_leaf_350_CLK _04263_ VGND VGND VPWR VPWR registers\[49\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21375_ _07309_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__buf_2
X_23114_ net64 VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__clkbuf_8
X_20326_ registers\[24\]\[55\] registers\[25\]\[55\] registers\[26\]\[55\] registers\[27\]\[55\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__mux4_1
X_24094_ _09634_ registers\[5\]\[57\] _10216_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__mux2_1
XFILLER_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28971_ registers\[24\]\[27\] _10361_ _12883_ VGND VGND VPWR VPWR _12891_ sky130_fd_sc_hd__mux2_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_289_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_289_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23045_ _09626_ registers\[62\]\[53\] _09620_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__mux2_1
X_27922_ _12339_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__clkbuf_1
X_20257_ _05069_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__buf_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27853_ registers\[32\]\[9\] _10323_ _12293_ VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__mux2_1
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ registers\[12\]\[51\] registers\[13\]\[51\] registers\[14\]\[51\] registers\[15\]\[51\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__mux4_1
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26804_ _11719_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkbuf_1
XTAP_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27784_ registers\[33\]\[40\] _10388_ _12266_ VGND VGND VPWR VPWR _12267_ sky130_fd_sc_hd__mux2_1
X_24996_ _10733_ registers\[52\]\[1\] _10731_ VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__mux2_1
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29523_ registers\[20\]\[1\] _12937_ _13211_ VGND VGND VPWR VPWR _13213_ sky130_fd_sc_hd__mux2_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26735_ _11683_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_1
X_23947_ _10146_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_801 _08973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_461_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_461_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_812 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29454_ _13176_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26666_ _11646_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_823 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23878_ _09554_ registers\[60\]\[19\] _10100_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__mux2_1
XFILLER_232_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_834 _09160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_845 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28405_ _12593_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__clkbuf_1
X_22829_ registers\[8\]\[62\] registers\[9\]\[62\] registers\[10\]\[62\] registers\[11\]\[62\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__mux4_1
XANTENNA_856 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25617_ _11093_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_867 _09364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29385_ _13139_ VGND VGND VPWR VPWR _13140_ sky130_fd_sc_hd__buf_4
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_878 _09529_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26597_ _11610_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_889 _09619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_213_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_213_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_198_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28336_ registers\[2\]\[46\] _10401_ _12550_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__mux2_1
X_16350_ _14531_ VGND VGND VPWR VPWR _14856_ sky130_fd_sc_hd__buf_4
XFILLER_242_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25548_ _11055_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16281_ _14528_ _14787_ _14788_ _14537_ VGND VGND VPWR VPWR _14789_ sky130_fd_sc_hd__a22o_1
X_25479_ _11019_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__clkbuf_1
X_28267_ registers\[2\]\[13\] _10332_ _12517_ VGND VGND VPWR VPWR _12521_ sky130_fd_sc_hd__mux2_1
XFILLER_185_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18020_ registers\[0\]\[55\] registers\[1\]\[55\] registers\[2\]\[55\] registers\[3\]\[55\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__mux4_1
XFILLER_185_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27218_ _11790_ registers\[37\]\[29\] _11958_ VGND VGND VPWR VPWR _11968_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28198_ _12484_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27149_ _11931_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30160_ _13547_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__clkbuf_1
X_19971_ registers\[12\]\[45\] registers\[13\]\[45\] registers\[14\]\[45\] registers\[15\]\[45\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__mux4_1
XFILLER_119_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18922_ _05666_ _05669_ _05508_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__o21ba_1
X_30091_ _13511_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1200 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1211 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1222 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18853_ registers\[28\]\[13\] registers\[29\]\[13\] registers\[30\]\[13\] registers\[31\]\[13\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__mux4_1
XANTENNA_1233 _00034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1244 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1255 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1266 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ registers\[48\]\[49\] registers\[49\]\[49\] registers\[50\]\[49\] registers\[51\]\[49\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__mux4_1
XTAP_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1277 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33850_ clknet_leaf_301_CLK _01964_ VGND VGND VPWR VPWR registers\[3\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_18784_ registers\[20\]\[11\] registers\[21\]\[11\] registers\[22\]\[11\] registers\[23\]\[11\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__mux4_1
XANTENNA_1288 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1299 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15996_ _14509_ VGND VGND VPWR VPWR _14510_ sky130_fd_sc_hd__buf_12
XTAP_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32801_ clknet_leaf_44_CLK _00915_ VGND VGND VPWR VPWR registers\[55\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_17735_ registers\[52\]\[47\] registers\[53\]\[47\] registers\[54\]\[47\] registers\[55\]\[47\]
+ _04476_ _04477_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__mux4_1
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33781_ clknet_leaf_344_CLK _01895_ VGND VGND VPWR VPWR registers\[40\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_30993_ registers\[10\]\[58\] _13056_ _13977_ VGND VGND VPWR VPWR _13986_ sky130_fd_sc_hd__mux2_1
X_35520_ clknet_leaf_236_CLK _03634_ VGND VGND VPWR VPWR registers\[13\]\[50\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_452_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_452_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_224_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32732_ clknet_leaf_50_CLK _00846_ VGND VGND VPWR VPWR registers\[56\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_17666_ _14502_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__buf_6
XFILLER_211_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19405_ registers\[0\]\[29\] registers\[1\]\[29\] registers\[2\]\[29\] registers\[3\]\[29\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__mux4_1
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35451_ clknet_leaf_304_CLK _03565_ VGND VGND VPWR VPWR registers\[14\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_16617_ registers\[16\]\[15\] registers\[17\]\[15\] registers\[18\]\[15\] registers\[19\]\[15\]
+ _14808_ _14809_ VGND VGND VPWR VPWR _15116_ sky130_fd_sc_hd__mux4_1
X_32663_ clknet_leaf_69_CLK _00777_ VGND VGND VPWR VPWR registers\[57\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_17597_ registers\[52\]\[43\] registers\[53\]\[43\] registers\[54\]\[43\] registers\[55\]\[43\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__mux4_1
XFILLER_23_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_204_CLK clknet_6_54__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_204_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34402_ clknet_leaf_473_CLK _02516_ VGND VGND VPWR VPWR registers\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19336_ registers\[4\]\[27\] registers\[5\]\[27\] registers\[6\]\[27\] registers\[7\]\[27\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__mux4_1
X_31614_ registers\[63\]\[32\] net26 _14310_ VGND VGND VPWR VPWR _14313_ sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16548_ _14801_ _15047_ _15048_ _14804_ VGND VGND VPWR VPWR _15049_ sky130_fd_sc_hd__a22o_1
X_35382_ clknet_leaf_320_CLK _03496_ VGND VGND VPWR VPWR registers\[15\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_32594_ clknet_leaf_71_CLK _00708_ VGND VGND VPWR VPWR registers\[58\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34333_ clknet_leaf_492_CLK _02447_ VGND VGND VPWR VPWR registers\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31545_ _09511_ _09940_ VGND VGND VPWR VPWR _14276_ sky130_fd_sc_hd__nor2_8
X_19267_ _05693_ _06003_ _06004_ _05696_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a22o_1
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16479_ _14978_ _14981_ _14945_ VGND VGND VPWR VPWR _14982_ sky130_fd_sc_hd__o21ba_1
X_18218_ registers\[44\]\[62\] registers\[45\]\[62\] registers\[46\]\[62\] registers\[47\]\[62\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__mux4_1
X_34264_ clknet_leaf_86_CLK _02378_ VGND VGND VPWR VPWR registers\[32\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_31476_ _14240_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__clkbuf_1
X_19198_ _05069_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__buf_4
X_36003_ clknet_leaf_445_CLK _04117_ VGND VGND VPWR VPWR registers\[63\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33215_ clknet_leaf_200_CLK _01329_ VGND VGND VPWR VPWR registers\[4\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_18149_ registers\[28\]\[59\] registers\[29\]\[59\] registers\[30\]\[59\] registers\[31\]\[59\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__mux4_1
XFILLER_191_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30427_ _13688_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__clkbuf_1
X_34195_ clknet_leaf_120_CLK _02309_ VGND VGND VPWR VPWR registers\[33\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33146_ clknet_leaf_285_CLK _01260_ VGND VGND VPWR VPWR registers\[50\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_21160_ registers\[32\]\[14\] registers\[33\]\[14\] registers\[34\]\[14\] registers\[35\]\[14\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__mux4_1
X_30358_ _13652_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__clkbuf_1
X_20111_ registers\[0\]\[49\] registers\[1\]\[49\] registers\[2\]\[49\] registers\[3\]\[49\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux4_1
XFILLER_171_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33077_ clknet_leaf_328_CLK _01191_ VGND VGND VPWR VPWR registers\[51\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_21091_ _07281_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__buf_4
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30289_ _13615_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__clkbuf_1
X_20042_ registers\[4\]\[47\] registers\[5\]\[47\] registers\[6\]\[47\] registers\[7\]\[47\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__mux4_1
X_32028_ clknet_leaf_49_CLK _00206_ VGND VGND VPWR VPWR registers\[62\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24850_ _09644_ registers\[54\]\[62\] _10586_ VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__mux2_1
XFILLER_74_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23801_ _09613_ registers\[29\]\[47\] _10061_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__mux2_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24781_ _09575_ registers\[54\]\[29\] _10609_ VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__mux2_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33979_ clknet_leaf_282_CLK _02093_ VGND VGND VPWR VPWR registers\[37\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_21993_ registers\[16\]\[37\] registers\[17\]\[37\] registers\[18\]\[37\] registers\[19\]\[37\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__mux4_1
XFILLER_39_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_443_CLK clknet_6_12__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_443_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26520_ _11513_ VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__buf_6
X_23732_ _09544_ registers\[29\]\[14\] _10028_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__mux2_1
XANTENNA_108 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35718_ clknet_leaf_155_CLK _03832_ VGND VGND VPWR VPWR registers\[10\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20944_ _07433_ _07633_ _07634_ _07438_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__a22o_1
XANTENNA_119 _00049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23663_ registers\[61\]\[47\] _09791_ _09987_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__mux2_1
X_26451_ _10766_ registers\[42\]\[17\] _11525_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__mux2_1
X_20875_ registers\[44\]\[6\] registers\[45\]\[6\] registers\[46\]\[6\] registers\[47\]\[6\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__mux4_1
X_35649_ clknet_leaf_240_CLK _03763_ VGND VGND VPWR VPWR registers\[11\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22614_ _09012_ _09256_ _09257_ _09018_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__a22o_1
X_25402_ _10806_ registers\[50\]\[36\] _10970_ VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__mux2_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26382_ _11496_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__clkbuf_1
X_29170_ registers\[23\]\[38\] _13014_ _12998_ VGND VGND VPWR VPWR _13015_ sky130_fd_sc_hd__mux2_1
XFILLER_35_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23594_ registers\[61\]\[14\] _09687_ _09954_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__mux2_1
XFILLER_74_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25333_ _10737_ registers\[50\]\[3\] _10937_ VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__mux2_1
X_28121_ _11746_ registers\[30\]\[8\] _12435_ VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__mux2_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22545_ _09187_ _09190_ _09083_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__o21ba_1
XFILLER_210_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25264_ _10804_ registers\[51\]\[35\] _10898_ VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__mux2_1
X_28052_ _12407_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22476_ _08812_ _09122_ _09123_ _08815_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__a22o_1
XFILLER_154_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27003_ _11851_ registers\[3\]\[58\] _11835_ VGND VGND VPWR VPWR _11852_ sky130_fd_sc_hd__mux2_1
X_24215_ _10232_ VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__buf_6
X_21427_ registers\[0\]\[21\] registers\[1\]\[21\] registers\[2\]\[21\] registers\[3\]\[21\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__mux4_1
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25195_ _10735_ registers\[51\]\[2\] _10865_ VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__mux2_1
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24146_ _09550_ registers\[58\]\[17\] _10244_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__mux2_1
XFILLER_108_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21358_ registers\[24\]\[19\] registers\[25\]\[19\] registers\[26\]\[19\] registers\[27\]\[19\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__mux4_1
X_20309_ registers\[36\]\[55\] registers\[37\]\[55\] registers\[38\]\[55\] registers\[39\]\[55\]
+ _06742_ _06743_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__mux4_1
X_24077_ _09617_ registers\[5\]\[49\] _10205_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__mux2_1
X_28954_ registers\[24\]\[19\] _10344_ _12872_ VGND VGND VPWR VPWR _12882_ sky130_fd_sc_hd__mux2_1
X_21289_ registers\[28\]\[17\] registers\[29\]\[17\] registers\[30\]\[17\] registers\[31\]\[17\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__mux4_1
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23028_ net43 VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__clkbuf_4
X_27905_ _12330_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__clkbuf_1
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28885_ _11834_ registers\[25\]\[50\] _12845_ VGND VGND VPWR VPWR _12846_ sky130_fd_sc_hd__mux2_1
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27836_ _12294_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__clkbuf_1
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27767_ registers\[33\]\[32\] _10372_ _12255_ VGND VGND VPWR VPWR _12258_ sky130_fd_sc_hd__mux2_1
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24979_ _09638_ registers\[53\]\[59\] _10713_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__mux2_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_434_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_434_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_29506_ _13203_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__clkbuf_1
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17520_ _15677_ _04304_ _04305_ _15682_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a22o_1
XFILLER_217_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26718_ _11674_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27698_ _09653_ _09707_ VGND VGND VPWR VPWR _12221_ sky130_fd_sc_hd__nor2_8
XFILLER_206_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_620 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_631 _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_642 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29437_ _13167_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__clkbuf_1
X_17451_ registers\[48\]\[39\] registers\[49\]\[39\] registers\[50\]\[39\] registers\[51\]\[39\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _15926_ sky130_fd_sc_hd__mux4_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_653 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26649_ _11637_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_664 _05365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_675 _05761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16402_ registers\[4\]\[9\] registers\[5\]\[9\] registers\[6\]\[9\] registers\[7\]\[9\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _14907_ sky130_fd_sc_hd__mux4_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_686 _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29368_ _09810_ registers\[22\]\[56\] _13124_ VGND VGND VPWR VPWR _13131_ sky130_fd_sc_hd__mux2_1
XANTENNA_697 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17382_ registers\[52\]\[37\] registers\[53\]\[37\] registers\[54\]\[37\] registers\[55\]\[37\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _15859_ sky130_fd_sc_hd__mux4_1
XFILLER_246_1392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19121_ _05747_ _05861_ _05862_ _05753_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__a22o_1
X_16333_ registers\[24\]\[7\] registers\[25\]\[7\] registers\[26\]\[7\] registers\[27\]\[7\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14840_ sky130_fd_sc_hd__mux4_1
X_28319_ registers\[2\]\[38\] _10384_ _12539_ VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__mux2_1
XFILLER_201_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29299_ _09730_ registers\[22\]\[23\] _13091_ VGND VGND VPWR VPWR _13095_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31330_ _14163_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__clkbuf_1
X_19052_ registers\[0\]\[19\] registers\[1\]\[19\] registers\[2\]\[19\] registers\[3\]\[19\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__mux4_1
XFILLER_185_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16264_ registers\[16\]\[5\] registers\[17\]\[5\] registers\[18\]\[5\] registers\[19\]\[5\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _14773_ sky130_fd_sc_hd__mux4_1
XFILLER_158_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18003_ _04750_ _04759_ _04766_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__or4_4
XFILLER_200_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31261_ registers\[8\]\[57\] net53 _14119_ VGND VGND VPWR VPWR _14127_ sky130_fd_sc_hd__mux2_1
X_16195_ _14570_ _14704_ _14705_ _14582_ VGND VGND VPWR VPWR _14706_ sky130_fd_sc_hd__a22o_1
XFILLER_142_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33000_ clknet_leaf_423_CLK _01114_ VGND VGND VPWR VPWR registers\[52\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_30212_ registers\[15\]\[8\] _12951_ _13566_ VGND VGND VPWR VPWR _13575_ sky130_fd_sc_hd__mux2_1
XFILLER_153_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31192_ registers\[8\]\[24\] net17 _14086_ VGND VGND VPWR VPWR _14091_ sky130_fd_sc_hd__mux2_1
XFILLER_113_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19954_ _06569_ _06670_ _06671_ _06574_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__a22o_1
X_30143_ _13538_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18905_ _05412_ _05651_ _05652_ _05416_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__a22o_1
X_34951_ clknet_leaf_208_CLK _03065_ VGND VGND VPWR VPWR registers\[22\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30074_ _13502_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__clkbuf_1
X_19885_ _06605_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_1030 _12934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1041 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1052 _13423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18836_ _05404_ _05584_ _05585_ _05410_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a22o_1
XANTENNA_1063 _13992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33902_ clknet_leaf_355_CLK _02016_ VGND VGND VPWR VPWR registers\[38\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34882_ clknet_leaf_229_CLK _02996_ VGND VGND VPWR VPWR registers\[23\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1074 _14418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1085 _14502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1096 _14524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33833_ clknet_leaf_458_CLK _01947_ VGND VGND VPWR VPWR registers\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_43__f_CLK clknet_5_21_0_CLK VGND VGND VPWR VPWR clknet_6_43__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_222_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18767_ registers\[48\]\[11\] registers\[49\]\[11\] registers\[50\]\[11\] registers\[51\]\[11\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux4_1
X_15979_ _14492_ VGND VGND VPWR VPWR _14493_ sky130_fd_sc_hd__buf_12
XFILLER_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_425_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_425_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_224_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17718_ _04294_ _04497_ _04498_ _04299_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__a22o_1
XFILLER_23_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33764_ clknet_leaf_56_CLK _01878_ VGND VGND VPWR VPWR registers\[40\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_30976_ _13921_ VGND VGND VPWR VPWR _13977_ sky130_fd_sc_hd__buf_4
X_18698_ registers\[8\]\[9\] registers\[9\]\[9\] registers\[10\]\[9\] registers\[11\]\[9\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__mux4_1
XFILLER_93_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_224_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32715_ clknet_leaf_165_CLK _00829_ VGND VGND VPWR VPWR registers\[57\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35503_ clknet_leaf_375_CLK _03617_ VGND VGND VPWR VPWR registers\[13\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_17649_ _04428_ _04431_ _04301_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__o21ba_1
XFILLER_23_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33695_ clknet_leaf_33_CLK _01809_ VGND VGND VPWR VPWR registers\[41\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35434_ clknet_leaf_398_CLK _03548_ VGND VGND VPWR VPWR registers\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_32646_ clknet_leaf_236_CLK _00760_ VGND VGND VPWR VPWR registers\[58\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20660_ _07358_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__buf_6
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19319_ registers\[44\]\[27\] registers\[45\]\[27\] registers\[46\]\[27\] registers\[47\]\[27\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__mux4_2
XFILLER_17_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35365_ clknet_leaf_462_CLK _03479_ VGND VGND VPWR VPWR registers\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_20591_ _07289_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__buf_4
X_32577_ clknet_leaf_233_CLK _00691_ VGND VGND VPWR VPWR registers\[5\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34316_ clknet_leaf_171_CLK _02430_ VGND VGND VPWR VPWR registers\[32\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_22330_ _08976_ _08981_ _08740_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__o21ba_1
X_31528_ _14267_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35296_ clknet_leaf_2_CLK _03410_ VGND VGND VPWR VPWR registers\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34247_ clknet_leaf_243_CLK _02361_ VGND VGND VPWR VPWR registers\[33\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22261_ _08669_ _08913_ _08914_ _08675_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__a22o_1
XFILLER_121_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31459_ _14231_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24000_ _09540_ registers\[5\]\[12\] _10172_ VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__mux2_1
X_21212_ registers\[12\]\[15\] registers\[13\]\[15\] registers\[14\]\[15\] registers\[15\]\[15\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__mux4_1
X_34178_ clknet_leaf_247_CLK _02292_ VGND VGND VPWR VPWR registers\[34\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22192_ _08844_ _08847_ _08740_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__o21ba_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21143_ _07581_ _07827_ _07828_ _07584_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__a22o_1
X_33129_ clknet_leaf_424_CLK _01243_ VGND VGND VPWR VPWR registers\[50\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25951_ _10806_ registers\[46\]\[36\] _11263_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__mux2_1
X_21074_ registers\[0\]\[11\] registers\[1\]\[11\] registers\[2\]\[11\] registers\[3\]\[11\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__mux4_1
XFILLER_101_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20025_ registers\[44\]\[47\] registers\[45\]\[47\] registers\[46\]\[47\] registers\[47\]\[47\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__mux4_1
X_24902_ _09561_ registers\[53\]\[22\] _10680_ VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28670_ _11755_ registers\[26\]\[12\] _12730_ VGND VGND VPWR VPWR _12733_ sky130_fd_sc_hd__mux2_1
X_25882_ _10737_ registers\[46\]\[3\] _11230_ VGND VGND VPWR VPWR _11234_ sky130_fd_sc_hd__mux2_1
XFILLER_189_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27621_ registers\[34\]\[27\] _10361_ _12173_ VGND VGND VPWR VPWR _12181_ sky130_fd_sc_hd__mux2_1
X_24833_ _10646_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_416_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_416_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27552_ _12143_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__clkbuf_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24764_ _10610_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__clkbuf_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _08469_ _08634_ _08637_ _08472_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__a22o_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1021 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26503_ _11560_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__clkbuf_1
X_20927_ registers\[0\]\[7\] registers\[1\]\[7\] registers\[2\]\[7\] registers\[3\]\[7\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__mux4_1
X_23715_ _09527_ registers\[29\]\[6\] _10017_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__mux2_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24695_ _09626_ registers\[55\]\[53\] _10569_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_0_0_CLK sky130_fd_sc_hd__clkbuf_8
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27483_ _12107_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__clkbuf_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29222_ net51 VGND VGND VPWR VPWR _13050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26434_ _10749_ registers\[42\]\[9\] _11514_ VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__mux2_1
XFILLER_159_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _07343_ _07550_ _07551_ _07353_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__a22o_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23646_ registers\[61\]\[39\] _09773_ _09976_ VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__mux2_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29153_ _13003_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__clkbuf_1
X_23577_ registers\[61\]\[6\] _09670_ _09943_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__mux2_1
XFILLER_70_1126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26365_ _10814_ registers\[43\]\[40\] _11487_ VGND VGND VPWR VPWR _11488_ sky130_fd_sc_hd__mux2_1
X_20789_ registers\[0\]\[3\] registers\[1\]\[3\] registers\[2\]\[3\] registers\[3\]\[3\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__mux4_1
XFILLER_122_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28104_ _12434_ VGND VGND VPWR VPWR _12435_ sky130_fd_sc_hd__buf_4
X_22528_ registers\[24\]\[52\] registers\[25\]\[52\] registers\[26\]\[52\] registers\[27\]\[52\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__mux4_1
XFILLER_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25316_ _10856_ registers\[51\]\[60\] _10864_ VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__mux2_1
X_26296_ _11451_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
X_29084_ registers\[23\]\[10\] _12955_ _12956_ VGND VGND VPWR VPWR _12957_ sky130_fd_sc_hd__mux2_1
XFILLER_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28035_ _11795_ registers\[31\]\[31\] _12397_ VGND VGND VPWR VPWR _12399_ sky130_fd_sc_hd__mux2_1
X_22459_ _09104_ _09105_ _09106_ _09107_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__a22o_1
XFILLER_183_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25247_ _10787_ registers\[51\]\[27\] _10887_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__mux2_1
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_902 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25178_ _10856_ registers\[52\]\[60\] _10730_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__mux2_1
XFILLER_108_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24129_ _09533_ registers\[58\]\[9\] _10233_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__mux2_1
X_29986_ registers\[17\]\[29\] _12995_ _13446_ VGND VGND VPWR VPWR _13456_ sky130_fd_sc_hd__mux2_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28937_ _12873_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16951_ _15341_ _15438_ _15439_ _15344_ VGND VGND VPWR VPWR _15440_ sky130_fd_sc_hd__a22o_1
XFILLER_89_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19670_ registers\[32\]\[37\] registers\[33\]\[37\] registers\[34\]\[37\] registers\[35\]\[37\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__mux4_1
XFILLER_81_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16882_ _15334_ _15371_ _15372_ _15339_ VGND VGND VPWR VPWR _15373_ sky130_fd_sc_hd__a22o_1
X_28868_ _11818_ registers\[25\]\[42\] _12834_ VGND VGND VPWR VPWR _12837_ sky130_fd_sc_hd__mux2_1
XFILLER_49_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18621_ _05077_ _05375_ _05376_ _05086_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__a22o_1
X_27819_ registers\[33\]\[57\] _10424_ _12277_ VGND VGND VPWR VPWR _12285_ sky130_fd_sc_hd__mux2_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28799_ _12800_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__clkbuf_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_407_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_407_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _05089_ _05308_ _05309_ _05100_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__a22o_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30830_ _13900_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ registers\[24\]\[40\] registers\[25\]\[40\] registers\[26\]\[40\] registers\[27\]\[40\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__mux4_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18483_ _05077_ _05241_ _05242_ _05086_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__a22o_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30761_ _13864_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_450 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32500_ clknet_leaf_353_CLK _00614_ VGND VGND VPWR VPWR registers\[60\]\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_461 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_472 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17434_ _15633_ _15908_ _15909_ _15636_ VGND VGND VPWR VPWR _15910_ sky130_fd_sc_hd__a22o_1
X_33480_ clknet_leaf_250_CLK _01594_ VGND VGND VPWR VPWR registers\[45\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_483 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30692_ registers\[12\]\[43\] _13025_ _13824_ VGND VGND VPWR VPWR _13828_ sky130_fd_sc_hd__mux2_1
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_494 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_221_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32431_ clknet_leaf_394_CLK _00545_ VGND VGND VPWR VPWR registers\[29\]\[33\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_19 _00029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17365_ _15638_ _15841_ _15842_ _15643_ VGND VGND VPWR VPWR _15843_ sky130_fd_sc_hd__a22o_1
XFILLER_53_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19104_ _05156_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__clkbuf_4
X_16316_ registers\[36\]\[7\] registers\[37\]\[7\] registers\[38\]\[7\] registers\[39\]\[7\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _14823_ sky130_fd_sc_hd__mux4_1
X_35150_ clknet_leaf_114_CLK _03264_ VGND VGND VPWR VPWR registers\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32362_ clknet_leaf_408_CLK _00476_ VGND VGND VPWR VPWR registers\[61\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17296_ _15772_ _15775_ _15645_ VGND VGND VPWR VPWR _15776_ sky130_fd_sc_hd__o21ba_1
XFILLER_105_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34101_ clknet_leaf_343_CLK _02215_ VGND VGND VPWR VPWR registers\[35\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31313_ _14154_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__clkbuf_1
X_19035_ registers\[40\]\[19\] registers\[41\]\[19\] registers\[42\]\[19\] registers\[43\]\[19\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__mux4_1
X_35081_ clknet_leaf_212_CLK _03195_ VGND VGND VPWR VPWR registers\[20\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16247_ registers\[56\]\[5\] registers\[57\]\[5\] registers\[58\]\[5\] registers\[59\]\[5\]
+ _14723_ _14532_ VGND VGND VPWR VPWR _14756_ sky130_fd_sc_hd__mux4_1
XFILLER_220_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32293_ clknet_leaf_446_CLK _00407_ VGND VGND VPWR VPWR registers\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_34032_ clknet_leaf_357_CLK _02146_ VGND VGND VPWR VPWR registers\[36\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_31244_ registers\[8\]\[49\] net44 _14108_ VGND VGND VPWR VPWR _14118_ sky130_fd_sc_hd__mux2_1
Xoutput104 net104 VGND VGND VPWR VPWR D1[22] sky130_fd_sc_hd__buf_2
X_16178_ registers\[36\]\[3\] registers\[37\]\[3\] registers\[38\]\[3\] registers\[39\]\[3\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14689_ sky130_fd_sc_hd__mux4_1
Xoutput115 net115 VGND VGND VPWR VPWR D1[32] sky130_fd_sc_hd__buf_2
XFILLER_173_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput126 net126 VGND VGND VPWR VPWR D1[42] sky130_fd_sc_hd__buf_2
XFILLER_86_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput137 net137 VGND VGND VPWR VPWR D1[52] sky130_fd_sc_hd__buf_2
Xoutput148 net148 VGND VGND VPWR VPWR D1[62] sky130_fd_sc_hd__buf_2
XFILLER_173_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput159 net159 VGND VGND VPWR VPWR D2[14] sky130_fd_sc_hd__buf_2
XFILLER_138_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31175_ registers\[8\]\[16\] net8 _14075_ VGND VGND VPWR VPWR _14082_ sky130_fd_sc_hd__mux2_1
XFILLER_82_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30126_ registers\[16\]\[31\] _13000_ _13528_ VGND VGND VPWR VPWR _13530_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19937_ registers\[12\]\[44\] registers\[13\]\[44\] registers\[14\]\[44\] registers\[15\]\[44\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__mux4_1
X_35983_ clknet_leaf_175_CLK _04097_ VGND VGND VPWR VPWR registers\[63\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30057_ registers\[17\]\[63\] _13066_ _13423_ VGND VGND VPWR VPWR _13493_ sky130_fd_sc_hd__mux2_1
X_34934_ clknet_leaf_307_CLK _03048_ VGND VGND VPWR VPWR registers\[22\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_19868_ registers\[8\]\[42\] registers\[9\]\[42\] registers\[10\]\[42\] registers\[11\]\[42\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__mux4_1
XFILLER_210_1019 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18819_ _05141_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__buf_6
X_34865_ clknet_leaf_385_CLK _02979_ VGND VGND VPWR VPWR registers\[23\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_19799_ _06379_ _06520_ _06521_ _06382_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__a22o_1
XFILLER_243_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21830_ _08491_ _08496_ _08430_ VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__o21ba_1
XFILLER_23_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33816_ clknet_leaf_11_CLK _01930_ VGND VGND VPWR VPWR registers\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_34796_ clknet_leaf_386_CLK _02910_ VGND VGND VPWR VPWR registers\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33747_ clknet_leaf_135_CLK _01861_ VGND VGND VPWR VPWR registers\[40\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_21761_ _07398_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__buf_2
X_30959_ _13968_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20712_ _07404_ _07409_ _07310_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__o21ba_1
X_23500_ _09908_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__clkbuf_1
X_24480_ _10458_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
X_33678_ clknet_leaf_147_CLK _01792_ VGND VGND VPWR VPWR registers\[41\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_21692_ _08119_ _08358_ _08361_ _08124_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__a22o_1
X_23431_ _09872_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20643_ _07323_ _07337_ _07339_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__o211a_1
X_35417_ clknet_leaf_14_CLK _03531_ VGND VGND VPWR VPWR registers\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_32629_ clknet_leaf_327_CLK _00743_ VGND VGND VPWR VPWR registers\[58\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26150_ _10735_ registers\[44\]\[2\] _11372_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__mux2_1
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35348_ clknet_leaf_79_CLK _03462_ VGND VGND VPWR VPWR registers\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_23362_ _09834_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
X_20574_ _07273_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22313_ _07317_ VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__buf_4
X_25101_ _10804_ registers\[52\]\[35\] _10794_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__mux2_1
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26081_ _11338_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
X_35279_ clknet_leaf_116_CLK _03393_ VGND VGND VPWR VPWR registers\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23293_ _09790_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25032_ net5 VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__buf_2
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22244_ registers\[16\]\[44\] registers\[17\]\[44\] registers\[18\]\[44\] registers\[19\]\[44\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__mux4_1
XFILLER_127_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29840_ _13379_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22175_ registers\[24\]\[42\] registers\[25\]\[42\] registers\[26\]\[42\] registers\[27\]\[42\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21126_ _07812_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
X_29771_ registers\[1\]\[55\] _13050_ _13337_ VGND VGND VPWR VPWR _13343_ sky130_fd_sc_hd__mux2_1
X_26983_ _11838_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1072 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28722_ _11807_ registers\[26\]\[37\] _12752_ VGND VGND VPWR VPWR _12760_ sky130_fd_sc_hd__mux2_1
XFILLER_87_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21057_ _07712_ _07721_ _07731_ _07745_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__or4_1
X_25934_ _10789_ registers\[46\]\[28\] _11252_ VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20008_ _05130_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__buf_4
X_28653_ _11738_ registers\[26\]\[4\] _12719_ VGND VGND VPWR VPWR _12724_ sky130_fd_sc_hd__mux2_1
XFILLER_59_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25865_ _11224_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27604_ registers\[34\]\[19\] _10344_ _12162_ VGND VGND VPWR VPWR _12172_ sky130_fd_sc_hd__mux2_1
X_24816_ _10637_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28584_ _12687_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25796_ _11188_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27535_ _11837_ registers\[35\]\[51\] _12133_ VGND VGND VPWR VPWR _12135_ sky130_fd_sc_hd__mux2_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24747_ _10601_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21959_ _07377_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__buf_6
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27466_ _12098_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24678_ _09609_ registers\[55\]\[45\] _10558_ VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__mux2_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29205_ _13038_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__clkbuf_1
X_26417_ _11515_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__clkbuf_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23629_ _09977_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27397_ _12006_ VGND VGND VPWR VPWR _12062_ sky130_fd_sc_hd__buf_4
XFILLER_74_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29136_ registers\[23\]\[27\] _12991_ _12977_ VGND VGND VPWR VPWR _12992_ sky130_fd_sc_hd__mux2_1
X_17150_ registers\[24\]\[30\] registers\[25\]\[30\] registers\[26\]\[30\] registers\[27\]\[30\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15634_ sky130_fd_sc_hd__mux4_1
X_26348_ _10798_ registers\[43\]\[32\] _11476_ VGND VGND VPWR VPWR _11479_ sky130_fd_sc_hd__mux2_1
Xinput17 DW[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_4
X_16101_ _14599_ _14612_ _14614_ VGND VGND VPWR VPWR _14615_ sky130_fd_sc_hd__o21ba_1
Xinput28 DW[34] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput39 DW[44] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_8
X_29067_ net56 VGND VGND VPWR VPWR _12945_ sky130_fd_sc_hd__buf_2
XFILLER_6_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17081_ _15290_ _15565_ _15566_ _15293_ VGND VGND VPWR VPWR _15567_ sky130_fd_sc_hd__a22o_1
Xclkbuf_6_7__f_CLK clknet_5_3_0_CLK VGND VGND VPWR VPWR clknet_6_7__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_26279_ _09868_ _11157_ VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__nand2_8
XFILLER_100_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16032_ _14492_ VGND VGND VPWR VPWR _14546_ sky130_fd_sc_hd__buf_12
X_28018_ _11778_ registers\[31\]\[23\] _12386_ VGND VGND VPWR VPWR _12390_ sky130_fd_sc_hd__mux2_1
XFILLER_164_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17983_ registers\[60\]\[54\] registers\[61\]\[54\] registers\[62\]\[54\] registers\[63\]\[54\]
+ _04755_ _04549_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__mux4_1
X_29969_ _13447_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__clkbuf_1
X_19722_ _06440_ _06446_ _06169_ _06170_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__o211a_1
X_16934_ _15420_ _15423_ _15288_ VGND VGND VPWR VPWR _15424_ sky130_fd_sc_hd__o21ba_1
X_32980_ clknet_leaf_64_CLK _01094_ VGND VGND VPWR VPWR registers\[52\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31931_ _14479_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__clkbuf_1
X_19653_ registers\[12\]\[36\] registers\[13\]\[36\] registers\[14\]\[36\] registers\[15\]\[36\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__mux4_1
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16865_ registers\[12\]\[22\] registers\[13\]\[22\] registers\[14\]\[22\] registers\[15\]\[22\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15357_ sky130_fd_sc_hd__mux4_1
XFILLER_238_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18604_ registers\[28\]\[6\] registers\[29\]\[6\] registers\[30\]\[6\] registers\[31\]\[6\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__mux4_1
X_34650_ clknet_leaf_20_CLK _02764_ VGND VGND VPWR VPWR registers\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_19584_ registers\[12\]\[34\] registers\[13\]\[34\] registers\[14\]\[34\] registers\[15\]\[34\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__mux4_1
X_31862_ _14443_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__clkbuf_1
X_16796_ _14587_ VGND VGND VPWR VPWR _15290_ sky130_fd_sc_hd__clkbuf_4
X_33601_ clknet_leaf_272_CLK _01715_ VGND VGND VPWR VPWR registers\[43\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18535_ registers\[20\]\[4\] registers\[21\]\[4\] registers\[22\]\[4\] registers\[23\]\[4\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__mux4_1
X_30813_ _13891_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34581_ clknet_leaf_95_CLK _02695_ VGND VGND VPWR VPWR registers\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31793_ registers\[59\]\[53\] net49 _14403_ VGND VGND VPWR VPWR _14407_ sky130_fd_sc_hd__mux2_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33532_ clknet_leaf_278_CLK _01646_ VGND VGND VPWR VPWR registers\[44\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_30744_ _13855_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__clkbuf_1
X_18466_ _05141_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__buf_6
XFILLER_179_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17417_ _14543_ VGND VGND VPWR VPWR _15893_ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33463_ clknet_leaf_340_CLK _01577_ VGND VGND VPWR VPWR registers\[45\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_18397_ _05159_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__buf_4
X_30675_ registers\[12\]\[35\] _13008_ _13813_ VGND VGND VPWR VPWR _13819_ sky130_fd_sc_hd__mux2_1
XFILLER_60_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35202_ clknet_leaf_222_CLK _03316_ VGND VGND VPWR VPWR registers\[18\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32414_ clknet_leaf_1_CLK _00528_ VGND VGND VPWR VPWR registers\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36182_ clknet_leaf_93_CLK _00126_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dfxtp_1
X_17348_ registers\[8\]\[36\] registers\[9\]\[36\] registers\[10\]\[36\] registers\[11\]\[36\]
+ _15792_ _15793_ VGND VGND VPWR VPWR _15826_ sky130_fd_sc_hd__mux4_1
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33394_ clknet_leaf_362_CLK _01508_ VGND VGND VPWR VPWR registers\[46\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35133_ clknet_leaf_299_CLK _03247_ VGND VGND VPWR VPWR registers\[1\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32345_ clknet_leaf_54_CLK _00459_ VGND VGND VPWR VPWR registers\[61\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17279_ _15549_ _15757_ _15758_ _15553_ VGND VGND VPWR VPWR _15759_ sky130_fd_sc_hd__a22o_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19018_ registers\[0\]\[18\] registers\[1\]\[18\] registers\[2\]\[18\] registers\[3\]\[18\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__mux4_1
X_35064_ clknet_leaf_309_CLK _03178_ VGND VGND VPWR VPWR registers\[20\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_20290_ registers\[12\]\[54\] registers\[13\]\[54\] registers\[14\]\[54\] registers\[15\]\[54\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__mux4_1
X_32276_ clknet_leaf_93_CLK _00390_ VGND VGND VPWR VPWR registers\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34015_ clknet_leaf_40_CLK _02129_ VGND VGND VPWR VPWR registers\[36\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_31227_ _14109_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_938 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31158_ registers\[8\]\[8\] net63 _14064_ VGND VGND VPWR VPWR _14073_ sky130_fd_sc_hd__mux2_1
XFILLER_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30109_ registers\[16\]\[23\] _12983_ _13517_ VGND VGND VPWR VPWR _13521_ sky130_fd_sc_hd__mux2_1
XFILLER_130_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23980_ _10164_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__clkbuf_1
X_35966_ clknet_leaf_197_CLK _04080_ VGND VGND VPWR VPWR registers\[6\]\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31089_ _14036_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34917_ clknet_leaf_447_CLK _03031_ VGND VGND VPWR VPWR registers\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_22931_ _09549_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
X_35897_ clknet_leaf_315_CLK _04011_ VGND VGND VPWR VPWR registers\[7\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_243_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25650_ registers\[48\]\[22\] _10351_ _11108_ VGND VGND VPWR VPWR _11111_ sky130_fd_sc_hd__mux2_1
X_22862_ registers\[12\]\[63\] registers\[13\]\[63\] registers\[14\]\[63\] registers\[15\]\[63\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__mux4_1
X_34848_ clknet_leaf_490_CLK _02962_ VGND VGND VPWR VPWR registers\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24601_ _10523_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21813_ _08334_ _08478_ _08479_ _08338_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__a22o_1
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25581_ registers\[4\]\[55\] _10420_ _11067_ VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__mux2_1
X_22793_ registers\[48\]\[61\] registers\[49\]\[61\] registers\[50\]\[61\] registers\[51\]\[61\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__mux4_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34779_ clknet_leaf_18_CLK _02893_ VGND VGND VPWR VPWR registers\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_212_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27320_ registers\[36\]\[13\] _10332_ _12018_ VGND VGND VPWR VPWR _12022_ sky130_fd_sc_hd__mux2_1
XFILLER_212_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21744_ registers\[12\]\[30\] registers\[13\]\[30\] registers\[14\]\[30\] registers\[15\]\[30\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__mux4_1
X_24532_ _09601_ registers\[56\]\[41\] _10484_ VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__mux2_1
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27251_ _11985_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__clkbuf_1
X_24463_ _10449_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
X_21675_ _07363_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__buf_4
XFILLER_237_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26202_ _10787_ registers\[44\]\[27\] _11394_ VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__mux2_1
X_23414_ _09861_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
X_20626_ _07324_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24394_ net43 VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__buf_4
X_27182_ _11949_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26133_ _11365_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
X_23345_ net60 VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__clkbuf_4
X_20557_ _05149_ _07255_ _07256_ _05159_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__a22o_1
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26064_ _11329_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
X_23276_ _09779_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
X_20488_ registers\[44\]\[61\] registers\[45\]\[61\] registers\[46\]\[61\] registers\[47\]\[61\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__mux4_1
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25015_ _10746_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
X_22227_ registers\[48\]\[44\] registers\[49\]\[44\] registers\[50\]\[44\] registers\[51\]\[44\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__mux4_1
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29823_ _13370_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__clkbuf_1
XTAP_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22158_ _07301_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_1607 _14581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1618 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1629 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21109_ registers\[8\]\[12\] registers\[9\]\[12\] registers\[10\]\[12\] registers\[11\]\[12\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__mux4_1
XTAP_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29754_ registers\[1\]\[47\] _13033_ _13326_ VGND VGND VPWR VPWR _13334_ sky130_fd_sc_hd__mux2_1
XFILLER_47_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22089_ _07338_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__clkbuf_4
X_26966_ _11826_ registers\[3\]\[46\] _11814_ VGND VGND VPWR VPWR _11827_ sky130_fd_sc_hd__mux2_1
XTAP_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28705_ _11790_ registers\[26\]\[29\] _12741_ VGND VGND VPWR VPWR _12751_ sky130_fd_sc_hd__mux2_1
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25917_ _11229_ VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__buf_4
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29685_ registers\[1\]\[14\] _12964_ _13293_ VGND VGND VPWR VPWR _13298_ sky130_fd_sc_hd__mux2_1
XFILLER_102_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26897_ net17 VGND VGND VPWR VPWR _11780_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28636_ _12714_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16650_ _15144_ _15145_ _15146_ _15147_ VGND VGND VPWR VPWR _15148_ sky130_fd_sc_hd__a22o_1
X_25848_ _10838_ registers\[47\]\[51\] _11214_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__mux2_1
XFILLER_47_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16581_ _15077_ _15080_ _14945_ VGND VGND VPWR VPWR _15081_ sky130_fd_sc_hd__o21ba_1
X_28567_ _12678_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25779_ _11179_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18320_ _05042_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__buf_4
X_27518_ _11820_ registers\[35\]\[43\] _12122_ VGND VGND VPWR VPWR _12126_ sky130_fd_sc_hd__mux2_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28498_ _11853_ registers\[28\]\[59\] _12632_ VGND VGND VPWR VPWR _12642_ sky130_fd_sc_hd__mux2_1
XFILLER_215_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_1187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _05011_ _05014_ _14524_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__o21ba_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27449_ _11750_ registers\[35\]\[10\] _12089_ VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__mux2_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17202_ _14539_ VGND VGND VPWR VPWR _15684_ sky130_fd_sc_hd__clkbuf_4
X_30460_ _13705_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__clkbuf_1
X_18182_ _04945_ _04948_ _14613_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__o21ba_1
XFILLER_54_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17133_ registers\[60\]\[30\] registers\[61\]\[30\] registers\[62\]\[30\] registers\[63\]\[30\]
+ _15413_ _15550_ VGND VGND VPWR VPWR _15617_ sky130_fd_sc_hd__mux4_1
X_29119_ _12980_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30391_ _13669_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32130_ clknet_leaf_461_CLK _00047_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17064_ _14543_ VGND VGND VPWR VPWR _15550_ sky130_fd_sc_hd__clkbuf_8
XFILLER_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16015_ _14492_ VGND VGND VPWR VPWR _14529_ sky130_fd_sc_hd__buf_12
X_32061_ clknet_leaf_288_CLK _00239_ VGND VGND VPWR VPWR registers\[62\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31012_ _13996_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35820_ clknet_leaf_391_CLK _03934_ VGND VGND VPWR VPWR registers\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_17966_ registers\[20\]\[53\] registers\[21\]\[53\] registers\[22\]\[53\] registers\[23\]\[53\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__mux4_1
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19705_ registers\[36\]\[38\] registers\[37\]\[38\] registers\[38\]\[38\] registers\[39\]\[38\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__mux4_1
X_16917_ _15341_ _15405_ _15406_ _15344_ VGND VGND VPWR VPWR _15407_ sky130_fd_sc_hd__a22o_1
X_32963_ clknet_leaf_266_CLK _01077_ VGND VGND VPWR VPWR registers\[53\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_35751_ clknet_leaf_459_CLK _03865_ VGND VGND VPWR VPWR registers\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17897_ _04637_ _04671_ _04672_ _04642_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__a22o_1
XFILLER_22_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_239_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34702_ clknet_leaf_111_CLK _02816_ VGND VGND VPWR VPWR registers\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31914_ _14470_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__clkbuf_1
X_19636_ _06233_ _06361_ _06362_ _06236_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__a22o_1
X_16848_ _15334_ _15337_ _15338_ _15339_ VGND VGND VPWR VPWR _15340_ sky130_fd_sc_hd__a22o_1
X_32894_ clknet_leaf_292_CLK _01008_ VGND VGND VPWR VPWR registers\[54\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_35682_ clknet_leaf_467_CLK _03796_ VGND VGND VPWR VPWR registers\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34633_ clknet_leaf_218_CLK _02747_ VGND VGND VPWR VPWR registers\[27\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31845_ _14434_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__clkbuf_1
X_19567_ _06226_ _06294_ _06295_ _06231_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__a22o_1
XFILLER_19_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16779_ _15198_ _15271_ _15272_ _15204_ VGND VGND VPWR VPWR _15273_ sky130_fd_sc_hd__a22o_1
XFILLER_230_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18518_ registers\[60\]\[4\] registers\[61\]\[4\] registers\[62\]\[4\] registers\[63\]\[4\]
+ _05276_ _05093_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__mux4_1
XFILLER_20_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34564_ clknet_leaf_206_CLK _02678_ VGND VGND VPWR VPWR registers\[28\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31776_ registers\[59\]\[45\] net40 _14392_ VGND VGND VPWR VPWR _14398_ sky130_fd_sc_hd__mux2_1
X_19498_ registers\[40\]\[32\] registers\[41\]\[32\] registers\[42\]\[32\] registers\[43\]\[32\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux4_1
XFILLER_90_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30727_ registers\[12\]\[60\] _13060_ _13779_ VGND VGND VPWR VPWR _13846_ sky130_fd_sc_hd__mux2_1
X_18449_ registers\[56\]\[2\] registers\[57\]\[2\] registers\[58\]\[2\] registers\[59\]\[2\]
+ _05079_ _05081_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__mux4_1
X_33515_ clknet_leaf_428_CLK _01629_ VGND VGND VPWR VPWR registers\[44\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_209_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34495_ clknet_leaf_296_CLK _02609_ VGND VGND VPWR VPWR registers\[2\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36234_ clknet_leaf_121_CLK _00120_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dfxtp_1
X_33446_ clknet_leaf_60_CLK _01560_ VGND VGND VPWR VPWR registers\[45\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_21460_ _07991_ _08135_ _08136_ _07995_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__a22o_1
XFILLER_147_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30658_ registers\[12\]\[27\] _12991_ _13802_ VGND VGND VPWR VPWR _13810_ sky130_fd_sc_hd__mux2_1
XFILLER_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20411_ _05040_ _07114_ _07115_ _05050_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__a22o_1
X_36165_ clknet_leaf_259_CLK _04279_ VGND VGND VPWR VPWR registers\[49\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_33377_ clknet_leaf_34_CLK _01491_ VGND VGND VPWR VPWR registers\[46\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_21391_ registers\[12\]\[20\] registers\[13\]\[20\] registers\[14\]\[20\] registers\[15\]\[20\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__mux4_1
X_30589_ _13773_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23130_ net6 VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__buf_6
X_32328_ clknet_leaf_153_CLK _00442_ VGND VGND VPWR VPWR registers\[19\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_20342_ registers\[56\]\[56\] registers\[57\]\[56\] registers\[58\]\[56\] registers\[59\]\[56\]
+ _06987_ _06777_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__mux4_1
X_35116_ clknet_leaf_388_CLK _03230_ VGND VGND VPWR VPWR registers\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36096_ clknet_leaf_267_CLK _04210_ VGND VGND VPWR VPWR registers\[59\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23061_ _09637_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
X_35047_ clknet_leaf_457_CLK _03161_ VGND VGND VPWR VPWR registers\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_20273_ _06912_ _06980_ _06981_ _06917_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__a22o_1
X_32259_ clknet_leaf_261_CLK _00373_ VGND VGND VPWR VPWR registers\[39\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_216_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22012_ _07328_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__clkbuf_4
XTAP_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_216_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26820_ _11727_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_1
XTAP_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26751_ registers\[40\]\[30\] _10367_ _11691_ VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__mux2_1
X_23963_ _10154_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35949_ clknet_leaf_392_CLK _04063_ VGND VGND VPWR VPWR registers\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25702_ registers\[48\]\[47\] _10403_ _11130_ VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29470_ _09775_ registers\[21\]\[40\] _13184_ VGND VGND VPWR VPWR _13185_ sky130_fd_sc_hd__mux2_1
X_22914_ net3 VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__buf_4
X_26682_ _11654_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23894_ _10118_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28421_ _11776_ registers\[28\]\[22\] _12599_ VGND VGND VPWR VPWR _12602_ sky130_fd_sc_hd__mux2_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25633_ registers\[48\]\[14\] _10334_ _11097_ VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__mux2_1
XFILLER_244_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22845_ registers\[40\]\[63\] registers\[41\]\[63\] registers\[42\]\[63\] registers\[43\]\[63\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__mux4_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_227_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28352_ _12565_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__clkbuf_1
X_25564_ registers\[4\]\[47\] _10403_ _11056_ VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__mux2_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22776_ registers\[24\]\[60\] registers\[25\]\[60\] registers\[26\]\[60\] registers\[27\]\[60\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__mux4_1
XFILLER_169_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27303_ registers\[36\]\[5\] _10315_ _12007_ VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__mux2_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24515_ _09584_ registers\[56\]\[33\] _10473_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28283_ _12529_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__clkbuf_1
X_21727_ _08126_ _08394_ _08395_ _08129_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__a22o_1
XFILLER_240_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25495_ registers\[4\]\[14\] _10334_ _11023_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__mux2_1
XFILLER_213_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27234_ _11976_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24446_ _09510_ registers\[56\]\[0\] _10440_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__mux2_1
X_21658_ _07326_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__buf_6
XFILLER_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20609_ _07296_ _07299_ _07302_ _07307_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__a22o_1
X_27165_ _11940_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24377_ registers\[57\]\[42\] _10393_ _10389_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__mux2_1
X_21589_ _07331_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__buf_6
XFILLER_201_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26116_ _10835_ registers\[45\]\[50\] _11356_ VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__mux2_1
X_23328_ registers\[9\]\[57\] _09813_ _09798_ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__mux2_1
XFILLER_165_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27096_ _11803_ registers\[38\]\[35\] _11898_ VGND VGND VPWR VPWR _11904_ sky130_fd_sc_hd__mux2_1
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26047_ _11320_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
X_23259_ registers\[39\]\[25\] _09742_ _09700_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1404 _00173_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1415 _00181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1426 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ registers\[28\]\[49\] registers\[29\]\[49\] registers\[30\]\[49\] registers\[31\]\[49\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__mux4_1
XTAP_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29806_ _13361_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1437 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1448 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27998_ _12379_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1459 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ _04527_ _04530_ _04301_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__o21ba_1
XFILLER_88_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26949_ _11815_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_1
X_29737_ registers\[1\]\[39\] _13016_ _13315_ VGND VGND VPWR VPWR _13325_ sky130_fd_sc_hd__mux2_1
XTAP_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16702_ _14527_ VGND VGND VPWR VPWR _15198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29668_ registers\[1\]\[6\] _12947_ _13282_ VGND VGND VPWR VPWR _13289_ sky130_fd_sc_hd__mux2_1
X_17682_ _04440_ _04447_ _04456_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__or4_2
XFILLER_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19421_ registers\[32\]\[30\] registers\[33\]\[30\] registers\[34\]\[30\] registers\[35\]\[30\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__mux4_1
X_28619_ _11839_ registers\[27\]\[52\] _12703_ VGND VGND VPWR VPWR _12706_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16633_ registers\[48\]\[16\] registers\[49\]\[16\] registers\[50\]\[16\] registers\[51\]\[16\]
+ _14858_ _14859_ VGND VGND VPWR VPWR _15131_ sky130_fd_sc_hd__mux4_1
XFILLER_169_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29599_ _13252_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31630_ _14276_ VGND VGND VPWR VPWR _14321_ sky130_fd_sc_hd__buf_4
XFILLER_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19352_ registers\[36\]\[28\] registers\[37\]\[28\] registers\[38\]\[28\] registers\[39\]\[28\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux4_1
XFILLER_216_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16564_ _14998_ _15062_ _15063_ _15001_ VGND VGND VPWR VPWR _15064_ sky130_fd_sc_hd__a22o_1
XFILLER_188_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18303_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__buf_4
XFILLER_200_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31561_ registers\[63\]\[7\] net62 _14277_ VGND VGND VPWR VPWR _14285_ sky130_fd_sc_hd__mux2_1
X_19283_ _05890_ _06018_ _06019_ _05893_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a22o_1
X_16495_ _14991_ _14994_ _14995_ _14996_ VGND VGND VPWR VPWR _14997_ sky130_fd_sc_hd__a22o_1
XFILLER_204_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33300_ clknet_leaf_125_CLK _01414_ VGND VGND VPWR VPWR registers\[47\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_18234_ _14511_ _04997_ _04998_ _14517_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a22o_1
X_30512_ _13733_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34280_ clknet_leaf_430_CLK _02394_ VGND VGND VPWR VPWR registers\[32\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31492_ _14248_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33231_ clknet_leaf_75_CLK _01345_ VGND VGND VPWR VPWR registers\[48\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_30443_ _09804_ registers\[14\]\[53\] _13693_ VGND VGND VPWR VPWR _13697_ sky130_fd_sc_hd__mux2_1
X_18165_ registers\[60\]\[60\] registers\[61\]\[60\] registers\[62\]\[60\] registers\[63\]\[60\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux4_1
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17116_ _15295_ _15599_ _15600_ _15300_ VGND VGND VPWR VPWR _15601_ sky130_fd_sc_hd__a22o_1
X_33162_ clknet_leaf_163_CLK _01276_ VGND VGND VPWR VPWR registers\[50\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_18096_ registers\[32\]\[58\] registers\[33\]\[58\] registers\[34\]\[58\] registers\[35\]\[58\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__mux4_1
XFILLER_209_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30374_ _09699_ registers\[14\]\[20\] _13660_ VGND VGND VPWR VPWR _13661_ sky130_fd_sc_hd__mux2_1
XFILLER_209_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32113_ clknet_leaf_467_CLK _00028_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17047_ _15533_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__clkbuf_1
X_33093_ clknet_leaf_258_CLK _01207_ VGND VGND VPWR VPWR registers\[51\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_32044_ clknet_leaf_374_CLK _00222_ VGND VGND VPWR VPWR registers\[62\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18998_ registers\[44\]\[18\] registers\[45\]\[18\] registers\[46\]\[18\] registers\[47\]\[18\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__mux4_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35803_ clknet_leaf_14_CLK _03917_ VGND VGND VPWR VPWR registers\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17949_ registers\[60\]\[53\] registers\[61\]\[53\] registers\[62\]\[53\] registers\[63\]\[53\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux4_1
XFILLER_117_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33995_ clknet_leaf_158_CLK _02109_ VGND VGND VPWR VPWR registers\[37\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35734_ clknet_leaf_87_CLK _03848_ VGND VGND VPWR VPWR registers\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_20960_ registers\[52\]\[8\] registers\[53\]\[8\] registers\[54\]\[8\] registers\[55\]\[8\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__mux4_1
XFILLER_187_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32946_ clknet_leaf_356_CLK _01060_ VGND VGND VPWR VPWR registers\[53\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19619_ registers\[4\]\[35\] registers\[5\]\[35\] registers\[6\]\[35\] registers\[7\]\[35\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__mux4_1
XFILLER_54_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35665_ clknet_leaf_109_CLK _03779_ VGND VGND VPWR VPWR registers\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_20891_ _07352_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__buf_4
XFILLER_241_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32877_ clknet_leaf_374_CLK _00991_ VGND VGND VPWR VPWR registers\[54\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_22630_ registers\[20\]\[55\] registers\[21\]\[55\] registers\[22\]\[55\] registers\[23\]\[55\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__mux4_1
XFILLER_198_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34616_ clknet_leaf_427_CLK _02730_ VGND VGND VPWR VPWR registers\[27\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_31828_ _14425_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__clkbuf_1
X_35596_ clknet_leaf_150_CLK _03710_ VGND VGND VPWR VPWR registers\[12\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22561_ _09201_ _09206_ _09102_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1043 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31759_ registers\[59\]\[37\] net31 _14381_ VGND VGND VPWR VPWR _14389_ sky130_fd_sc_hd__mux2_1
X_34547_ clknet_leaf_414_CLK _02661_ VGND VGND VPWR VPWR registers\[28\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24300_ _10341_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
X_21512_ registers\[40\]\[24\] registers\[41\]\[24\] registers\[42\]\[24\] registers\[43\]\[24\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__mux4_1
XFILLER_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22492_ registers\[24\]\[51\] registers\[25\]\[51\] registers\[26\]\[51\] registers\[27\]\[51\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__mux4_1
X_25280_ _10912_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34478_ clknet_leaf_389_CLK _02592_ VGND VGND VPWR VPWR registers\[2\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24231_ _10296_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
X_36217_ clknet_leaf_115_CLK _00101_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dfxtp_1
X_21443_ _07278_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__clkbuf_8
X_33429_ clknet_leaf_123_CLK _01543_ VGND VGND VPWR VPWR registers\[45\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24162_ _10260_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
X_36148_ clknet_leaf_350_CLK _04262_ VGND VGND VPWR VPWR registers\[49\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_21374_ _07783_ _08051_ _08052_ _07786_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__a22o_1
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23113_ _09675_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
X_20325_ _07029_ _07032_ _06866_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__o21ba_1
X_24093_ _10223_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
X_28970_ _12890_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36079_ clknet_leaf_371_CLK _04193_ VGND VGND VPWR VPWR registers\[59\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23044_ net49 VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__buf_4
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27921_ registers\[32\]\[41\] _10391_ _12337_ VGND VGND VPWR VPWR _12339_ sky130_fd_sc_hd__mux2_1
X_20256_ _05067_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__buf_6
XFILLER_162_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_755 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27852_ _12302_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ _06717_ _06897_ _06898_ _06720_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__a22o_1
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26803_ registers\[40\]\[55\] _10420_ _11713_ VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__mux2_1
XTAP_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27783_ _12221_ VGND VGND VPWR VPWR _12266_ sky130_fd_sc_hd__buf_4
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24995_ net12 VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_29_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29522_ _13212_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__clkbuf_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26734_ registers\[40\]\[22\] _10351_ _11680_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__mux2_1
X_23946_ _09622_ registers\[60\]\[51\] _10144_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__mux2_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_802 _08973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29453_ _09758_ registers\[21\]\[32\] _13173_ VGND VGND VPWR VPWR _13176_ sky130_fd_sc_hd__mux2_1
Xclkbuf_5_6_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_6_0_CLK sky130_fd_sc_hd__clkbuf_8
X_26665_ _10844_ registers\[41\]\[54\] _11641_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__mux2_1
XFILLER_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_813 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_824 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ _10109_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_835 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28404_ _11759_ registers\[28\]\[14\] _12588_ VGND VGND VPWR VPWR _12593_ sky130_fd_sc_hd__mux2_1
XFILLER_233_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_846 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25616_ registers\[48\]\[6\] _10317_ _11086_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__mux2_1
XANTENNA_857 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29384_ _09866_ _10015_ VGND VGND VPWR VPWR _13139_ sky130_fd_sc_hd__nand2_8
X_22828_ _09461_ _09464_ _07338_ _07340_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__o211a_1
XFILLER_44_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_868 _09364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26596_ _10775_ registers\[41\]\[21\] _11608_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__mux2_1
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_879 _09538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28335_ _12556_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25547_ registers\[4\]\[39\] _10386_ _11045_ VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22759_ registers\[36\]\[60\] registers\[37\]\[60\] registers\[38\]\[60\] registers\[39\]\[60\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__mux4_1
XFILLER_125_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16280_ registers\[48\]\[6\] registers\[49\]\[6\] registers\[50\]\[6\] registers\[51\]\[6\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _14788_ sky130_fd_sc_hd__mux4_1
X_28266_ _12520_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__clkbuf_1
X_25478_ registers\[4\]\[6\] _10317_ _11012_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27217_ _11967_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__clkbuf_1
X_24429_ registers\[57\]\[59\] _10428_ _10410_ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28197_ _11822_ registers\[30\]\[44\] _12479_ VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__mux2_1
XFILLER_139_985 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27148_ _11855_ registers\[38\]\[60\] _11864_ VGND VGND VPWR VPWR _11931_ sky130_fd_sc_hd__mux2_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1001 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19970_ _06374_ _06686_ _06687_ _06377_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a22o_1
XFILLER_126_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27079_ _11786_ registers\[38\]\[27\] _11887_ VGND VGND VPWR VPWR _11895_ sky130_fd_sc_hd__mux2_1
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18921_ _05501_ _05667_ _05668_ _05506_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__a22o_1
XTAP_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30090_ registers\[16\]\[14\] _12964_ _13506_ VGND VGND VPWR VPWR _13511_ sky130_fd_sc_hd__mux2_1
XFILLER_79_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1201 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1212 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1223 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1234 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18852_ _05496_ _05600_ _05601_ _05499_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__a22o_1
XFILLER_84_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1245 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1256 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17803_ registers\[56\]\[49\] registers\[57\]\[49\] registers\[58\]\[49\] registers\[59\]\[49\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__mux4_1
XFILLER_132_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1267 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1278 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18783_ registers\[28\]\[11\] registers\[29\]\[11\] registers\[30\]\[11\] registers\[31\]\[11\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__mux4_1
XFILLER_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _14508_ VGND VGND VPWR VPWR _14509_ sky130_fd_sc_hd__buf_2
XANTENNA_1289 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ registers\[60\]\[47\] registers\[61\]\[47\] registers\[62\]\[47\] registers\[63\]\[47\]
+ _04412_ _15893_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__mux4_1
X_32800_ clknet_leaf_44_CLK _00914_ VGND VGND VPWR VPWR registers\[55\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30992_ _13985_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__clkbuf_1
X_33780_ clknet_leaf_346_CLK _01894_ VGND VGND VPWR VPWR registers\[40\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_247_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17665_ _04443_ _04446_ _15963_ _15964_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__o211a_1
X_32731_ clknet_leaf_52_CLK _00845_ VGND VGND VPWR VPWR registers\[56\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19404_ registers\[8\]\[29\] registers\[9\]\[29\] registers\[10\]\[29\] registers\[11\]\[29\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__mux4_1
X_16616_ registers\[24\]\[15\] registers\[25\]\[15\] registers\[26\]\[15\] registers\[27\]\[15\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15115_ sky130_fd_sc_hd__mux4_1
X_32662_ clknet_leaf_69_CLK _00776_ VGND VGND VPWR VPWR registers\[57\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35450_ clknet_leaf_304_CLK _03564_ VGND VGND VPWR VPWR registers\[14\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_986 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17596_ registers\[60\]\[43\] registers\[61\]\[43\] registers\[62\]\[43\] registers\[63\]\[43\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__mux4_1
XFILLER_108_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34401_ clknet_leaf_488_CLK _02515_ VGND VGND VPWR VPWR registers\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_31613_ _14312_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19335_ registers\[12\]\[27\] registers\[13\]\[27\] registers\[14\]\[27\] registers\[15\]\[27\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__mux4_1
X_16547_ registers\[4\]\[13\] registers\[5\]\[13\] registers\[6\]\[13\] registers\[7\]\[13\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15048_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32593_ clknet_leaf_73_CLK _00707_ VGND VGND VPWR VPWR registers\[58\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_35381_ clknet_leaf_323_CLK _03495_ VGND VGND VPWR VPWR registers\[15\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31544_ _14275_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__clkbuf_1
X_19266_ registers\[4\]\[25\] registers\[5\]\[25\] registers\[6\]\[25\] registers\[7\]\[25\]
+ _05766_ _05767_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__mux4_1
X_34332_ clknet_leaf_0_CLK _02446_ VGND VGND VPWR VPWR registers\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_16478_ _14801_ _14979_ _14980_ _14804_ VGND VGND VPWR VPWR _14981_ sky130_fd_sc_hd__a22o_1
X_18217_ _14528_ _04980_ _04981_ _14537_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__a22o_1
X_34263_ clknet_leaf_106_CLK _02377_ VGND VGND VPWR VPWR registers\[32\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31475_ _09753_ registers\[6\]\[30\] _14239_ VGND VGND VPWR VPWR _14240_ sky130_fd_sc_hd__mux2_1
X_19197_ _05067_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__buf_4
X_33214_ clknet_leaf_198_CLK _01328_ VGND VGND VPWR VPWR registers\[4\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_36002_ clknet_leaf_444_CLK _04116_ VGND VGND VPWR VPWR registers\[63\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_18148_ _04632_ _04914_ _04915_ _04635_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__a22o_1
XFILLER_145_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30426_ _09786_ registers\[14\]\[45\] _13682_ VGND VGND VPWR VPWR _13688_ sky130_fd_sc_hd__mux2_1
X_34194_ clknet_leaf_122_CLK _02308_ VGND VGND VPWR VPWR registers\[33\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33145_ clknet_leaf_285_CLK _01259_ VGND VGND VPWR VPWR registers\[50\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_18079_ registers\[8\]\[57\] registers\[9\]\[57\] registers\[10\]\[57\] registers\[11\]\[57\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__mux4_1
X_30357_ _09683_ registers\[14\]\[12\] _13649_ VGND VGND VPWR VPWR _13652_ sky130_fd_sc_hd__mux2_1
XFILLER_105_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20110_ registers\[8\]\[49\] registers\[9\]\[49\] registers\[10\]\[49\] registers\[11\]\[49\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__mux4_1
XFILLER_131_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33076_ clknet_leaf_350_CLK _01190_ VGND VGND VPWR VPWR registers\[51\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_21090_ _07278_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__buf_4
X_30288_ registers\[15\]\[44\] _13027_ _13610_ VGND VGND VPWR VPWR _13615_ sky130_fd_sc_hd__mux2_1
XFILLER_113_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20041_ registers\[12\]\[47\] registers\[13\]\[47\] registers\[14\]\[47\] registers\[15\]\[47\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__mux4_1
X_32027_ clknet_leaf_54_CLK _00205_ VGND VGND VPWR VPWR registers\[62\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_140_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_140_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1790 _14584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23800_ _10068_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24780_ _10618_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
X_33978_ clknet_leaf_281_CLK _02092_ VGND VGND VPWR VPWR registers\[37\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_21992_ registers\[24\]\[37\] registers\[25\]\[37\] registers\[26\]\[37\] registers\[27\]\[37\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__mux4_1
XFILLER_82_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35717_ clknet_leaf_216_CLK _03831_ VGND VGND VPWR VPWR registers\[10\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23731_ _10032_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ registers\[32\]\[8\] registers\[33\]\[8\] registers\[34\]\[8\] registers\[35\]\[8\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__mux4_1
XFILLER_226_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_109 _00048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32929_ clknet_leaf_44_CLK _01043_ VGND VGND VPWR VPWR registers\[53\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26450_ _11532_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__clkbuf_1
X_35648_ clknet_leaf_244_CLK _03762_ VGND VGND VPWR VPWR registers\[11\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23662_ _09994_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _07433_ _07565_ _07566_ _07438_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__a22o_1
XFILLER_198_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25401_ _10976_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__clkbuf_1
X_22613_ registers\[48\]\[55\] registers\[49\]\[55\] registers\[50\]\[55\] registers\[51\]\[55\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__mux4_1
X_26381_ _10831_ registers\[43\]\[48\] _11487_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__mux2_1
XFILLER_197_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35579_ clknet_leaf_305_CLK _03693_ VGND VGND VPWR VPWR registers\[12\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_23593_ _09958_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_1
X_28120_ _12443_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25332_ _10940_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__clkbuf_1
X_22544_ _09155_ _09188_ _09189_ _09158_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__a22o_1
XFILLER_14_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28051_ _11811_ registers\[31\]\[39\] _12397_ VGND VGND VPWR VPWR _12407_ sky130_fd_sc_hd__mux2_1
X_25263_ _10903_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__clkbuf_1
X_22475_ registers\[36\]\[51\] registers\[37\]\[51\] registers\[38\]\[51\] registers\[39\]\[51\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__mux4_1
XFILLER_241_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27002_ net54 VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24214_ _10287_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
X_21426_ registers\[8\]\[21\] registers\[9\]\[21\] registers\[10\]\[21\] registers\[11\]\[21\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__mux4_1
X_25194_ _10867_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21357_ _08033_ _08036_ _07730_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__o21ba_1
X_24145_ _10251_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20308_ registers\[44\]\[55\] registers\[45\]\[55\] registers\[46\]\[55\] registers\[47\]\[55\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__mux4_1
X_24076_ _10214_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__clkbuf_1
X_21288_ _07732_ _07968_ _07969_ _07735_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__a22o_1
X_28953_ _12881_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__clkbuf_1
X_20239_ registers\[40\]\[53\] registers\[41\]\[53\] registers\[42\]\[53\] registers\[43\]\[53\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__mux4_1
X_23027_ _09614_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27904_ registers\[32\]\[33\] _10374_ _12326_ VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__mux2_1
X_28884_ _12789_ VGND VGND VPWR VPWR _12845_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_131_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_131_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27835_ registers\[32\]\[0\] _10303_ _12293_ VGND VGND VPWR VPWR _12294_ sky130_fd_sc_hd__mux2_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27766_ _12257_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__clkbuf_1
X_24978_ _10722_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__clkbuf_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29505_ _09813_ registers\[21\]\[57\] _13195_ VGND VGND VPWR VPWR _13203_ sky130_fd_sc_hd__mux2_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26717_ registers\[40\]\[14\] _10334_ _11669_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__mux2_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _09605_ registers\[60\]\[43\] _10133_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__mux2_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27697_ _12220_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__clkbuf_1
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_610 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_621 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29436_ _09740_ registers\[21\]\[24\] _13162_ VGND VGND VPWR VPWR _13167_ sky130_fd_sc_hd__mux2_1
XANTENNA_632 _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17450_ registers\[56\]\[39\] registers\[57\]\[39\] registers\[58\]\[39\] registers\[59\]\[39\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _15925_ sky130_fd_sc_hd__mux4_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_643 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26648_ _10827_ registers\[41\]\[46\] _11630_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__mux2_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_654 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_665 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16401_ registers\[12\]\[9\] registers\[13\]\[9\] registers\[14\]\[9\] registers\[15\]\[9\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14906_ sky130_fd_sc_hd__mux4_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_676 _05794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29367_ _13130_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_687 _06292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17381_ registers\[60\]\[37\] registers\[61\]\[37\] registers\[62\]\[37\] registers\[63\]\[37\]
+ _15756_ _15550_ VGND VGND VPWR VPWR _15858_ sky130_fd_sc_hd__mux4_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_198_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_198_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26579_ _10758_ registers\[41\]\[13\] _11597_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__mux2_1
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_698 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19120_ registers\[48\]\[21\] registers\[49\]\[21\] registers\[50\]\[21\] registers\[51\]\[21\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__mux4_1
X_16332_ _14835_ _14838_ _14585_ VGND VGND VPWR VPWR _14839_ sky130_fd_sc_hd__o21ba_1
X_28318_ _12547_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29298_ _13094_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19051_ registers\[8\]\[19\] registers\[9\]\[19\] registers\[10\]\[19\] registers\[11\]\[19\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__mux4_1
XFILLER_51_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28249_ _12511_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__clkbuf_1
X_16263_ registers\[24\]\[5\] registers\[25\]\[5\] registers\[26\]\[5\] registers\[27\]\[5\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14772_ sky130_fd_sc_hd__mux4_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18002_ _04771_ _04774_ _04644_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__o21ba_1
X_31260_ _14126_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16194_ registers\[4\]\[3\] registers\[5\]\[3\] registers\[6\]\[3\] registers\[7\]\[3\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14705_ sky130_fd_sc_hd__mux4_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30211_ _13574_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31191_ _14090_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_370_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_370_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30142_ registers\[16\]\[39\] _13016_ _13528_ VGND VGND VPWR VPWR _13538_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19953_ registers\[32\]\[45\] registers\[33\]\[45\] registers\[34\]\[45\] registers\[35\]\[45\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__mux4_1
XFILLER_206_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18904_ registers\[52\]\[15\] registers\[53\]\[15\] registers\[54\]\[15\] registers\[55\]\[15\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__mux4_1
XFILLER_45_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_122_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34950_ clknet_leaf_208_CLK _03064_ VGND VGND VPWR VPWR registers\[22\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_30073_ registers\[16\]\[6\] _12947_ _13495_ VGND VGND VPWR VPWR _13502_ sky130_fd_sc_hd__mux2_1
X_19884_ _06581_ _06588_ _06595_ _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__or4_4
XFILLER_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1020 _12434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1031 _12934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1042 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1053 _13494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33901_ clknet_leaf_325_CLK _02015_ VGND VGND VPWR VPWR registers\[38\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18835_ registers\[48\]\[13\] registers\[49\]\[13\] registers\[50\]\[13\] registers\[51\]\[13\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__mux4_1
XTAP_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34881_ clknet_leaf_203_CLK _02995_ VGND VGND VPWR VPWR registers\[23\]\[51\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1064 _14063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1075 _14474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1086 _14502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1097 _14527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33832_ clknet_leaf_457_CLK _01946_ VGND VGND VPWR VPWR registers\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15978_ net65 VGND VGND VPWR VPWR _14492_ sky130_fd_sc_hd__buf_8
X_18766_ registers\[56\]\[11\] registers\[57\]\[11\] registers\[58\]\[11\] registers\[59\]\[11\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__mux4_1
XFILLER_114_1471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17717_ registers\[20\]\[46\] registers\[21\]\[46\] registers\[22\]\[46\] registers\[23\]\[46\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__mux4_1
X_30975_ _13976_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__clkbuf_1
X_33763_ clknet_leaf_48_CLK _01877_ VGND VGND VPWR VPWR registers\[40\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_18697_ _05447_ _05450_ _05103_ _05105_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__o211a_1
X_35502_ clknet_leaf_393_CLK _03616_ VGND VGND VPWR VPWR registers\[13\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32714_ clknet_leaf_161_CLK _00828_ VGND VGND VPWR VPWR registers\[57\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_17648_ _04294_ _04429_ _04430_ _04299_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__a22o_1
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33694_ clknet_leaf_27_CLK _01808_ VGND VGND VPWR VPWR registers\[41\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35433_ clknet_leaf_398_CLK _03547_ VGND VGND VPWR VPWR registers\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_32645_ clknet_leaf_264_CLK _00759_ VGND VGND VPWR VPWR registers\[58\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_17579_ _14578_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_189_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_189_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19318_ _05883_ _06052_ _06053_ _05888_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a22o_1
X_20590_ _07280_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__buf_12
X_32576_ clknet_leaf_231_CLK _00690_ VGND VGND VPWR VPWR registers\[5\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35364_ clknet_leaf_467_CLK _03478_ VGND VGND VPWR VPWR registers\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_866 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34315_ clknet_leaf_158_CLK _02429_ VGND VGND VPWR VPWR registers\[32\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_31527_ _09808_ registers\[6\]\[55\] _14261_ VGND VGND VPWR VPWR _14267_ sky130_fd_sc_hd__mux2_1
X_19249_ registers\[44\]\[25\] registers\[45\]\[25\] registers\[46\]\[25\] registers\[47\]\[25\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__mux4_1
X_35295_ clknet_leaf_2_CLK _03409_ VGND VGND VPWR VPWR registers\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22260_ registers\[48\]\[45\] registers\[49\]\[45\] registers\[50\]\[45\] registers\[51\]\[45\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__mux4_1
XFILLER_30_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34246_ clknet_leaf_248_CLK _02360_ VGND VGND VPWR VPWR registers\[33\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_31458_ _09717_ registers\[6\]\[22\] _14228_ VGND VGND VPWR VPWR _14231_ sky130_fd_sc_hd__mux2_1
XFILLER_118_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21211_ _07581_ _07893_ _07894_ _07584_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__a22o_1
X_30409_ _09769_ registers\[14\]\[37\] _13671_ VGND VGND VPWR VPWR _13679_ sky130_fd_sc_hd__mux2_1
X_34177_ clknet_leaf_258_CLK _02291_ VGND VGND VPWR VPWR registers\[34\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_22191_ _08812_ _08845_ _08846_ _08815_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__a22o_1
X_31389_ _14194_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_361_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_361_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21142_ registers\[0\]\[13\] registers\[1\]\[13\] registers\[2\]\[13\] registers\[3\]\[13\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__mux4_1
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33128_ clknet_leaf_435_CLK _01242_ VGND VGND VPWR VPWR registers\[50\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_113_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25950_ _11269_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_21073_ registers\[8\]\[11\] registers\[9\]\[11\] registers\[10\]\[11\] registers\[11\]\[11\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__mux4_1
X_33059_ clknet_leaf_47_CLK _01173_ VGND VGND VPWR VPWR registers\[51\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20024_ _06569_ _06738_ _06739_ _06574_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__a22o_1
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24901_ _10682_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25881_ _11233_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
X_27620_ _12180_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24832_ _09626_ registers\[54\]\[53\] _10642_ VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__mux2_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27551_ _11853_ registers\[35\]\[59\] _12133_ VGND VGND VPWR VPWR _12143_ sky130_fd_sc_hd__mux2_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24763_ _09556_ registers\[54\]\[20\] _10609_ VGND VGND VPWR VPWR _10610_ sky130_fd_sc_hd__mux2_1
XFILLER_215_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ registers\[36\]\[37\] registers\[37\]\[37\] registers\[38\]\[37\] registers\[39\]\[37\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__mux4_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26502_ _10817_ registers\[42\]\[41\] _11558_ VGND VGND VPWR VPWR _11560_ sky130_fd_sc_hd__mux2_1
X_23714_ _10023_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20926_ registers\[8\]\[7\] registers\[9\]\[7\] registers\[10\]\[7\] registers\[11\]\[7\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__mux4_1
XFILLER_148_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27482_ _11784_ registers\[35\]\[26\] _12100_ VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__mux2_1
X_24694_ _10572_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29221_ _13049_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__clkbuf_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26433_ _11523_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_202_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _09985_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20857_ registers\[0\]\[5\] registers\[1\]\[5\] registers\[2\]\[5\] registers\[3\]\[5\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__mux4_1
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29152_ registers\[23\]\[32\] _13002_ _12998_ VGND VGND VPWR VPWR _13003_ sky130_fd_sc_hd__mux2_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26364_ _11442_ VGND VGND VPWR VPWR _11487_ sky130_fd_sc_hd__buf_4
X_23576_ _09949_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20788_ registers\[8\]\[3\] registers\[9\]\[3\] registers\[10\]\[3\] registers\[11\]\[3\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__mux4_1
X_28103_ _10014_ _10585_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__nand2_8
XFILLER_161_1255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25315_ _10930_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22527_ _09170_ _09173_ _09102_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__o21ba_1
X_29083_ _12934_ VGND VGND VPWR VPWR _12956_ sky130_fd_sc_hd__buf_4
X_26295_ _10745_ registers\[43\]\[7\] _11443_ VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__mux2_1
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28034_ _12398_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__clkbuf_1
X_25246_ _10894_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_1
X_22458_ _07352_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21409_ _08079_ _08086_ _08087_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__o21ba_1
X_25177_ net57 VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__buf_2
XFILLER_194_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_352_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_352_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22389_ registers\[20\]\[48\] registers\[21\]\[48\] registers\[22\]\[48\] registers\[23\]\[48\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__mux4_1
XFILLER_124_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24128_ _10242_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29985_ _13455_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_104_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28936_ registers\[24\]\[10\] _10325_ _12872_ VGND VGND VPWR VPWR _12873_ sky130_fd_sc_hd__mux2_1
X_16950_ registers\[36\]\[25\] registers\[37\]\[25\] registers\[38\]\[25\] registers\[39\]\[25\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15439_ sky130_fd_sc_hd__mux4_1
X_24059_ _09598_ registers\[5\]\[40\] _10205_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__mux2_1
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16881_ registers\[32\]\[23\] registers\[33\]\[23\] registers\[34\]\[23\] registers\[35\]\[23\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15372_ sky130_fd_sc_hd__mux4_1
X_28867_ _12836_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18620_ registers\[48\]\[7\] registers\[49\]\[7\] registers\[50\]\[7\] registers\[51\]\[7\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__mux4_1
X_27818_ _12284_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__clkbuf_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28798_ _11748_ registers\[25\]\[9\] _12790_ VGND VGND VPWR VPWR _12800_ sky130_fd_sc_hd__mux2_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ registers\[52\]\[5\] registers\[53\]\[5\] registers\[54\]\[5\] registers\[55\]\[5\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__mux4_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27749_ _12248_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__clkbuf_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17502_ _14490_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__buf_4
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ registers\[48\]\[3\] registers\[49\]\[3\] registers\[50\]\[3\] registers\[51\]\[3\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__mux4_1
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30760_ _09681_ registers\[11\]\[11\] _13862_ VGND VGND VPWR VPWR _13864_ sky130_fd_sc_hd__mux2_1
XFILLER_46_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_440 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_451 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ registers\[16\]\[38\] registers\[17\]\[38\] registers\[18\]\[38\] registers\[19\]\[38\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _15909_ sky130_fd_sc_hd__mux4_1
XANTENNA_462 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29419_ _09691_ registers\[21\]\[16\] _13151_ VGND VGND VPWR VPWR _13158_ sky130_fd_sc_hd__mux2_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_473 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30691_ _13827_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_484 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_495 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32430_ clknet_leaf_394_CLK _00544_ VGND VGND VPWR VPWR registers\[29\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17364_ registers\[20\]\[36\] registers\[21\]\[36\] registers\[22\]\[36\] registers\[23\]\[36\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15842_ sky130_fd_sc_hd__mux4_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_1396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16315_ _14573_ VGND VGND VPWR VPWR _14822_ sky130_fd_sc_hd__buf_6
X_19103_ _05079_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__buf_4
XFILLER_201_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32361_ clknet_leaf_452_CLK _00475_ VGND VGND VPWR VPWR registers\[61\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17295_ _15638_ _15773_ _15774_ _15643_ VGND VGND VPWR VPWR _15775_ sky130_fd_sc_hd__a22o_1
X_31312_ registers\[7\]\[17\] net9 _14146_ VGND VGND VPWR VPWR _14154_ sky130_fd_sc_hd__mux2_1
X_19034_ _05778_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
X_34100_ clknet_leaf_349_CLK _02214_ VGND VGND VPWR VPWR registers\[35\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_16246_ _14751_ _14754_ _14525_ VGND VGND VPWR VPWR _14755_ sky130_fd_sc_hd__o21ba_1
X_35080_ clknet_leaf_210_CLK _03194_ VGND VGND VPWR VPWR registers\[20\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32292_ clknet_leaf_446_CLK _00406_ VGND VGND VPWR VPWR registers\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34031_ clknet_leaf_357_CLK _02145_ VGND VGND VPWR VPWR registers\[36\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31243_ _14117_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__clkbuf_1
X_16177_ registers\[44\]\[3\] registers\[45\]\[3\] registers\[46\]\[3\] registers\[47\]\[3\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14688_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_343_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_343_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput105 net105 VGND VGND VPWR VPWR D1[23] sky130_fd_sc_hd__buf_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput116 net116 VGND VGND VPWR VPWR D1[33] sky130_fd_sc_hd__buf_2
Xoutput127 net127 VGND VGND VPWR VPWR D1[43] sky130_fd_sc_hd__buf_2
Xoutput138 net138 VGND VGND VPWR VPWR D1[53] sky130_fd_sc_hd__buf_2
XFILLER_177_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31174_ _14081_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__clkbuf_1
Xoutput149 net149 VGND VGND VPWR VPWR D1[63] sky130_fd_sc_hd__buf_2
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30125_ _13529_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__clkbuf_1
X_19936_ _06374_ _06653_ _06654_ _06377_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__a22o_1
X_35982_ clknet_leaf_178_CLK _04096_ VGND VGND VPWR VPWR registers\[63\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30056_ _13492_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34933_ clknet_leaf_384_CLK _03047_ VGND VGND VPWR VPWR registers\[22\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_19867_ _06584_ _06587_ _06512_ _06513_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__o211a_1
XFILLER_68_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18818_ _05496_ _05567_ _05568_ _05499_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__a22o_1
XFILLER_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34864_ clknet_leaf_388_CLK _02978_ VGND VGND VPWR VPWR registers\[23\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_19798_ registers\[4\]\[40\] registers\[5\]\[40\] registers\[6\]\[40\] registers\[7\]\[40\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__mux4_1
XFILLER_231_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33815_ clknet_leaf_88_CLK _01929_ VGND VGND VPWR VPWR registers\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18749_ registers\[28\]\[10\] registers\[29\]\[10\] registers\[30\]\[10\] registers\[31\]\[10\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__mux4_1
XFILLER_243_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34795_ clknet_leaf_451_CLK _02909_ VGND VGND VPWR VPWR registers\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33746_ clknet_leaf_128_CLK _01860_ VGND VGND VPWR VPWR registers\[40\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_21760_ _08423_ _08424_ _08427_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__a22o_1
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30958_ registers\[10\]\[41\] _13021_ _13966_ VGND VGND VPWR VPWR _13968_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20711_ _07296_ _07405_ _07408_ _07302_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__a22o_1
XFILLER_149_1386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33677_ clknet_leaf_76_CLK _01791_ VGND VGND VPWR VPWR registers\[42\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_21691_ registers\[32\]\[29\] registers\[33\]\[29\] registers\[34\]\[29\] registers\[35\]\[29\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__mux4_1
XFILLER_145_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30889_ _13931_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23430_ _09517_ registers\[19\]\[1\] _09870_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__mux2_1
X_35416_ clknet_leaf_13_CLK _03530_ VGND VGND VPWR VPWR registers\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_20642_ _07340_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__buf_2
XFILLER_71_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32628_ clknet_leaf_351_CLK _00742_ VGND VGND VPWR VPWR registers\[58\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20573_ _07251_ _07258_ _07265_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__or4_2
X_35347_ clknet_leaf_77_CLK _03461_ VGND VGND VPWR VPWR registers\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_23361_ registers\[39\]\[34\] _09762_ _09829_ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32559_ clknet_leaf_373_CLK _00673_ VGND VGND VPWR VPWR registers\[5\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_25100_ net29 VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__buf_2
XFILLER_176_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22312_ _07377_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__buf_6
X_26080_ _10800_ registers\[45\]\[33\] _11334_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__mux2_1
X_35278_ clknet_leaf_116_CLK _03392_ VGND VGND VPWR VPWR registers\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23292_ registers\[39\]\[26\] _09744_ _09700_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25031_ _10757_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22243_ registers\[24\]\[44\] registers\[25\]\[44\] registers\[26\]\[44\] registers\[27\]\[44\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__mux4_1
X_34229_ clknet_leaf_343_CLK _02343_ VGND VGND VPWR VPWR registers\[33\]\[39\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_334_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_334_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22174_ _08827_ _08830_ _08759_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21125_ _07788_ _07795_ _07802_ _07811_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__or4_2
X_29770_ _13342_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__clkbuf_1
X_26982_ _11837_ registers\[3\]\[51\] _11835_ VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__mux2_1
XFILLER_28_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25933_ _11260_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
X_28721_ _12759_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21056_ _07736_ _07743_ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__o21ba_1
XFILLER_87_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20007_ registers\[4\]\[46\] registers\[5\]\[46\] registers\[6\]\[46\] registers\[7\]\[46\]
+ _06452_ _06453_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__mux4_1
X_28652_ _12723_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25864_ _10854_ registers\[47\]\[59\] _11214_ VGND VGND VPWR VPWR _11224_ sky130_fd_sc_hd__mux2_1
XFILLER_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24815_ _09609_ registers\[54\]\[45\] _10631_ VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__mux2_1
X_27603_ _12171_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28583_ _11803_ registers\[27\]\[35\] _12681_ VGND VGND VPWR VPWR _12687_ sky130_fd_sc_hd__mux2_1
X_25795_ _10785_ registers\[47\]\[26\] _11181_ VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__mux2_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27534_ _12134_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__clkbuf_1
X_24746_ _09540_ registers\[54\]\[12\] _10598_ VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__mux2_1
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ registers\[24\]\[36\] registers\[25\]\[36\] registers\[26\]\[36\] registers\[27\]\[36\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__mux4_1
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20909_ _07601_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27465_ _11767_ registers\[35\]\[18\] _12089_ VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__mux2_1
XFILLER_163_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24677_ _10563_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21889_ _07349_ VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__buf_4
XFILLER_202_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26416_ _10728_ registers\[42\]\[0\] _11514_ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__mux2_1
XFILLER_159_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29204_ registers\[23\]\[49\] _13037_ _13019_ VGND VGND VPWR VPWR _13038_ sky130_fd_sc_hd__mux2_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23628_ registers\[61\]\[30\] _09753_ _09976_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__mux2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27396_ _12061_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29135_ net20 VGND VGND VPWR VPWR _12991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26347_ _11478_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__clkbuf_1
X_23559_ _09646_ registers\[19\]\[63\] _09869_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16100_ _14613_ VGND VGND VPWR VPWR _14614_ sky130_fd_sc_hd__clkbuf_4
Xinput18 DW[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
XFILLER_195_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29066_ _12944_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput29 DW[35] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
X_17080_ registers\[16\]\[28\] registers\[17\]\[28\] registers\[18\]\[28\] registers\[19\]\[28\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15566_ sky130_fd_sc_hd__mux4_1
X_26278_ _11441_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16031_ registers\[60\]\[0\] registers\[61\]\[0\] registers\[62\]\[0\] registers\[63\]\[0\]
+ _14542_ _14544_ VGND VGND VPWR VPWR _14545_ sky130_fd_sc_hd__mux4_1
X_28017_ _12389_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25229_ _10885_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_325_CLK clknet_6_44__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_325_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17982_ _14541_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__buf_6
X_29968_ registers\[17\]\[20\] _12976_ _13446_ VGND VGND VPWR VPWR _13447_ sky130_fd_sc_hd__mux2_1
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19721_ _06441_ _06443_ _06444_ _06445_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__a22o_1
XFILLER_81_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28919_ registers\[24\]\[2\] _10309_ _12861_ VGND VGND VPWR VPWR _12864_ sky130_fd_sc_hd__mux2_1
XFILLER_172_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16933_ _15144_ _15421_ _15422_ _15147_ VGND VGND VPWR VPWR _15423_ sky130_fd_sc_hd__a22o_1
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29899_ _13410_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31930_ _09806_ registers\[49\]\[54\] _14474_ VGND VGND VPWR VPWR _14479_ sky130_fd_sc_hd__mux2_1
X_19652_ _05059_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__buf_4
X_16864_ _15139_ _15354_ _15355_ _15142_ VGND VGND VPWR VPWR _15356_ sky130_fd_sc_hd__a22o_1
XFILLER_237_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18603_ _05137_ _05356_ _05359_ _05147_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a22o_1
XFILLER_225_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16795_ _15284_ _15287_ _15288_ VGND VGND VPWR VPWR _15289_ sky130_fd_sc_hd__o21ba_1
X_19583_ _06031_ _06310_ _06311_ _06034_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__a22o_1
X_31861_ _09702_ registers\[49\]\[21\] _14441_ VGND VGND VPWR VPWR _14443_ sky130_fd_sc_hd__mux2_1
XFILLER_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33600_ clknet_leaf_272_CLK _01714_ VGND VGND VPWR VPWR registers\[43\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18534_ registers\[28\]\[4\] registers\[29\]\[4\] registers\[30\]\[4\] registers\[31\]\[4\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__mux4_1
X_30812_ _09766_ registers\[11\]\[36\] _13884_ VGND VGND VPWR VPWR _13891_ sky130_fd_sc_hd__mux2_1
X_31792_ _14406_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__clkbuf_1
X_34580_ clknet_leaf_94_CLK _02694_ VGND VGND VPWR VPWR registers\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33531_ clknet_leaf_279_CLK _01645_ VGND VGND VPWR VPWR registers\[44\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_18465_ _05137_ _05224_ _05225_ _05147_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a22o_1
X_30743_ _09664_ registers\[11\]\[3\] _13851_ VGND VGND VPWR VPWR _13855_ sky130_fd_sc_hd__mux2_1
XANTENNA_270 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_1428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_292 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17416_ _14539_ VGND VGND VPWR VPWR _15892_ sky130_fd_sc_hd__clkbuf_4
X_18396_ _05064_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__buf_12
X_30674_ _13818_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__clkbuf_1
X_33462_ clknet_leaf_341_CLK _01576_ VGND VGND VPWR VPWR registers\[45\]\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35201_ clknet_leaf_221_CLK _03315_ VGND VGND VPWR VPWR registers\[18\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32413_ clknet_leaf_492_CLK _00527_ VGND VGND VPWR VPWR registers\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17347_ _14490_ VGND VGND VPWR VPWR _15825_ sky130_fd_sc_hd__buf_4
XFILLER_174_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36181_ clknet_leaf_93_CLK _00125_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33393_ clknet_leaf_361_CLK _01507_ VGND VGND VPWR VPWR registers\[46\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35132_ clknet_leaf_299_CLK _03246_ VGND VGND VPWR VPWR registers\[1\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32344_ clknet_leaf_54_CLK _00458_ VGND VGND VPWR VPWR registers\[61\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_17278_ registers\[52\]\[34\] registers\[53\]\[34\] registers\[54\]\[34\] registers\[55\]\[34\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15758_ sky130_fd_sc_hd__mux4_1
XFILLER_140_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16229_ _14562_ VGND VGND VPWR VPWR _14739_ sky130_fd_sc_hd__buf_6
X_19017_ registers\[8\]\[18\] registers\[9\]\[18\] registers\[10\]\[18\] registers\[11\]\[18\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__mux4_1
X_32275_ clknet_leaf_105_CLK _00389_ VGND VGND VPWR VPWR registers\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35063_ clknet_leaf_304_CLK _03177_ VGND VGND VPWR VPWR registers\[20\]\[41\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_316_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_316_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34014_ clknet_leaf_23_CLK _02128_ VGND VGND VPWR VPWR registers\[36\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31226_ registers\[8\]\[40\] net35 _14108_ VGND VGND VPWR VPWR _14109_ sky130_fd_sc_hd__mux2_1
XFILLER_142_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31157_ _14072_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30108_ _13520_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__clkbuf_1
X_19919_ registers\[32\]\[44\] registers\[33\]\[44\] registers\[34\]\[44\] registers\[35\]\[44\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__mux4_1
X_35965_ clknet_leaf_305_CLK _04079_ VGND VGND VPWR VPWR registers\[6\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31088_ registers\[0\]\[39\] _13016_ _14026_ VGND VGND VPWR VPWR _14036_ sky130_fd_sc_hd__mux2_1
XFILLER_69_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30039_ registers\[17\]\[54\] _13048_ _13479_ VGND VGND VPWR VPWR _13484_ sky130_fd_sc_hd__mux2_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34916_ clknet_leaf_473_CLK _03030_ VGND VGND VPWR VPWR registers\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_22930_ _09548_ registers\[62\]\[16\] _09536_ VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__mux2_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35896_ clknet_leaf_314_CLK _04010_ VGND VGND VPWR VPWR registers\[7\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22861_ _07276_ _09495_ _09496_ _07286_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__a22o_1
XFILLER_186_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34847_ clknet_leaf_488_CLK _02961_ VGND VGND VPWR VPWR registers\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24600_ _09531_ registers\[55\]\[8\] _10514_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__mux2_1
X_21812_ registers\[52\]\[32\] registers\[53\]\[32\] registers\[54\]\[32\] registers\[55\]\[32\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__mux4_1
X_25580_ _11072_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
X_22792_ registers\[56\]\[61\] registers\[57\]\[61\] registers\[58\]\[61\] registers\[59\]\[61\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__mux4_1
XFILLER_25_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34778_ clknet_leaf_19_CLK _02892_ VGND VGND VPWR VPWR registers\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_243_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_231_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24531_ _10485_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33729_ clknet_leaf_257_CLK _01843_ VGND VGND VPWR VPWR registers\[41\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21743_ _08267_ _08408_ _08411_ _08270_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__a22o_1
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27250_ _11822_ registers\[37\]\[44\] _11980_ VGND VGND VPWR VPWR _11985_ sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24462_ _09531_ registers\[56\]\[8\] _10440_ VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__mux2_1
XFILLER_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21674_ _07361_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__buf_6
XFILLER_40_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26201_ _11401_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23413_ registers\[39\]\[59\] _09817_ _09851_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__mux2_1
X_20625_ _07294_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__buf_12
X_27181_ _11753_ registers\[37\]\[11\] _11947_ VGND VGND VPWR VPWR _11949_ sky130_fd_sc_hd__mux2_1
X_24393_ _10404_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26132_ _10852_ registers\[45\]\[58\] _11356_ VGND VGND VPWR VPWR _11365_ sky130_fd_sc_hd__mux2_1
XFILLER_137_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23344_ _09824_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20556_ registers\[52\]\[63\] registers\[53\]\[63\] registers\[54\]\[63\] registers\[55\]\[63\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__mux4_1
X_26063_ _10783_ registers\[45\]\[25\] _11323_ VGND VGND VPWR VPWR _11329_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_307_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_307_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23275_ registers\[9\]\[41\] _09778_ _09776_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__mux2_1
X_20487_ _06912_ _07187_ _07188_ _06917_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__a22o_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25014_ _10745_ registers\[52\]\[7\] _10731_ VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22226_ registers\[56\]\[44\] registers\[57\]\[44\] registers\[58\]\[44\] registers\[59\]\[44\]
+ _08880_ _08670_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__mux4_1
XFILLER_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29822_ registers\[18\]\[15\] _12966_ _13364_ VGND VGND VPWR VPWR _13370_ sky130_fd_sc_hd__mux2_1
XTAP_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22157_ registers\[36\]\[42\] registers\[37\]\[42\] registers\[38\]\[42\] registers\[39\]\[42\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__mux4_1
XANTENNA_1608 _14581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1619 _15647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21108_ _07791_ _07794_ _07719_ _07720_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__o211a_1
XFILLER_121_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29753_ _13333_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26965_ net41 VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__clkbuf_4
X_22088_ _08677_ _08745_ _08746_ _08681_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__a22o_1
XTAP_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28704_ _12750_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25916_ _11251_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
X_21039_ registers\[4\]\[10\] registers\[5\]\[10\] registers\[6\]\[10\] registers\[7\]\[10\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__mux4_1
XFILLER_247_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29684_ _13297_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__clkbuf_1
X_26896_ _11779_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28635_ _11855_ registers\[27\]\[60\] _12647_ VGND VGND VPWR VPWR _12714_ sky130_fd_sc_hd__mux2_1
X_25847_ _11215_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16580_ _14801_ _15078_ _15079_ _14804_ VGND VGND VPWR VPWR _15080_ sky130_fd_sc_hd__a22o_1
XFILLER_216_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25778_ _10768_ registers\[47\]\[18\] _11170_ VGND VGND VPWR VPWR _11179_ sky130_fd_sc_hd__mux2_1
X_28566_ _11786_ registers\[27\]\[27\] _12670_ VGND VGND VPWR VPWR _12678_ sky130_fd_sc_hd__mux2_1
XFILLER_222_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24729_ _09523_ registers\[54\]\[4\] _10587_ VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__mux2_1
X_27517_ _12125_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__clkbuf_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28497_ _12641_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__clkbuf_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18250_ _14540_ _05012_ _05013_ _14551_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a22o_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27448_ _12077_ VGND VGND VPWR VPWR _12089_ sky130_fd_sc_hd__buf_6
XFILLER_54_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _15677_ _15680_ _15681_ _15682_ VGND VGND VPWR VPWR _15683_ sky130_fd_sc_hd__a22o_1
XFILLER_141_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18181_ _14570_ _04946_ _04947_ _14582_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__a22o_1
X_27379_ registers\[36\]\[41\] _10391_ _12051_ VGND VGND VPWR VPWR _12053_ sky130_fd_sc_hd__mux2_1
XFILLER_180_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17132_ _15541_ _15614_ _15615_ _15547_ VGND VGND VPWR VPWR _15616_ sky130_fd_sc_hd__a22o_1
XFILLER_8_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29118_ registers\[23\]\[21\] _12979_ _12977_ VGND VGND VPWR VPWR _12980_ sky130_fd_sc_hd__mux2_1
X_30390_ _09749_ registers\[14\]\[28\] _13660_ VGND VGND VPWR VPWR _13669_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29049_ _09651_ _09650_ _09649_ VGND VGND VPWR VPWR _12932_ sky130_fd_sc_hd__or3b_1
X_17063_ _14539_ VGND VGND VPWR VPWR _15549_ sky130_fd_sc_hd__buf_4
X_16014_ _14527_ VGND VGND VPWR VPWR _14528_ sky130_fd_sc_hd__buf_2
X_32060_ clknet_leaf_288_CLK _00238_ VGND VGND VPWR VPWR registers\[62\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31011_ registers\[0\]\[2\] _12939_ _13993_ VGND VGND VPWR VPWR _13996_ sky130_fd_sc_hd__mux2_1
XFILLER_174_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ registers\[28\]\[53\] registers\[29\]\[53\] registers\[30\]\[53\] registers\[31\]\[53\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__mux4_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19704_ registers\[44\]\[38\] registers\[45\]\[38\] registers\[46\]\[38\] registers\[47\]\[38\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux4_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35750_ clknet_leaf_463_CLK _03864_ VGND VGND VPWR VPWR registers\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16916_ registers\[36\]\[24\] registers\[37\]\[24\] registers\[38\]\[24\] registers\[39\]\[24\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15406_ sky130_fd_sc_hd__mux4_1
X_32962_ clknet_leaf_266_CLK _01076_ VGND VGND VPWR VPWR registers\[53\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17896_ registers\[20\]\[51\] registers\[21\]\[51\] registers\[22\]\[51\] registers\[23\]\[51\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__mux4_1
XFILLER_66_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34701_ clknet_leaf_148_CLK _02815_ VGND VGND VPWR VPWR registers\[26\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_31913_ _09788_ registers\[49\]\[46\] _14463_ VGND VGND VPWR VPWR _14470_ sky130_fd_sc_hd__mux2_1
X_19635_ registers\[36\]\[36\] registers\[37\]\[36\] registers\[38\]\[36\] registers\[39\]\[36\]
+ _06056_ _06057_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux4_1
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35681_ clknet_leaf_489_CLK _03795_ VGND VGND VPWR VPWR registers\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_16847_ _14500_ VGND VGND VPWR VPWR _15339_ sky130_fd_sc_hd__clkbuf_4
X_32893_ clknet_leaf_288_CLK _01007_ VGND VGND VPWR VPWR registers\[54\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34632_ clknet_leaf_218_CLK _02746_ VGND VGND VPWR VPWR registers\[27\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_241_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31844_ _09685_ registers\[49\]\[13\] _14430_ VGND VGND VPWR VPWR _14434_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19566_ registers\[32\]\[34\] registers\[33\]\[34\] registers\[34\]\[34\] registers\[35\]\[34\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16778_ registers\[48\]\[20\] registers\[49\]\[20\] registers\[50\]\[20\] registers\[51\]\[20\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15272_ sky130_fd_sc_hd__mux4_1
XFILLER_225_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18517_ _05090_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__buf_6
XFILLER_34_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34563_ clknet_leaf_205_CLK _02677_ VGND VGND VPWR VPWR registers\[28\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31775_ _14397_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__clkbuf_1
X_19497_ _05045_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__clkbuf_4
XFILLER_240_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33514_ clknet_leaf_428_CLK _01628_ VGND VGND VPWR VPWR registers\[44\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18448_ _05203_ _05208_ _05074_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__o21ba_1
X_30726_ _13845_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34494_ clknet_leaf_297_CLK _02608_ VGND VGND VPWR VPWR registers\[2\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36233_ clknet_leaf_121_CLK _00118_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dfxtp_1
X_33445_ clknet_leaf_59_CLK _01559_ VGND VGND VPWR VPWR registers\[45\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18379_ _05141_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__buf_6
X_30657_ _13809_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_93_CLK clknet_6_16__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_93_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20410_ registers\[0\]\[58\] registers\[1\]\[58\] registers\[2\]\[58\] registers\[3\]\[58\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__mux4_1
XFILLER_159_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36164_ clknet_leaf_260_CLK _04278_ VGND VGND VPWR VPWR registers\[49\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21390_ _07924_ _08065_ _08068_ _07927_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__a22o_1
X_30588_ _09815_ registers\[13\]\[58\] _13764_ VGND VGND VPWR VPWR _13773_ sky130_fd_sc_hd__mux2_1
XFILLER_119_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33376_ clknet_leaf_33_CLK _01490_ VGND VGND VPWR VPWR registers\[46\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35115_ clknet_leaf_459_CLK _03229_ VGND VGND VPWR VPWR registers\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32327_ clknet_leaf_153_CLK _00441_ VGND VGND VPWR VPWR registers\[19\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_20341_ _07044_ _07047_ _06847_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__o21ba_2
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36095_ clknet_leaf_290_CLK _04209_ VGND VGND VPWR VPWR registers\[59\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20272_ registers\[32\]\[54\] registers\[33\]\[54\] registers\[34\]\[54\] registers\[35\]\[54\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__mux4_1
XFILLER_190_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23060_ _09636_ registers\[62\]\[58\] _09620_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__mux2_1
X_35046_ clknet_leaf_456_CLK _03160_ VGND VGND VPWR VPWR registers\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32258_ clknet_leaf_261_CLK _00372_ VGND VGND VPWR VPWR registers\[39\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22011_ _07326_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__buf_4
XTAP_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31209_ registers\[8\]\[32\] net26 _14097_ VGND VGND VPWR VPWR _14100_ sky130_fd_sc_hd__mux2_1
X_32189_ clknet_leaf_465_CLK _00303_ VGND VGND VPWR VPWR registers\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26750_ _11657_ VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__buf_4
XFILLER_99_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23962_ _09638_ registers\[60\]\[59\] _10144_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__mux2_1
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35948_ clknet_leaf_394_CLK _04062_ VGND VGND VPWR VPWR registers\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_233_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25701_ _11137_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
X_22913_ _09537_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26681_ _10860_ registers\[41\]\[62\] _11585_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__mux2_1
X_35879_ clknet_leaf_457_CLK _03993_ VGND VGND VPWR VPWR registers\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_23893_ _09569_ registers\[60\]\[26\] _10111_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__mux2_1
XFILLER_216_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25632_ _11101_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
X_28420_ _12601_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22844_ _09480_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28351_ registers\[2\]\[53\] _10416_ _12561_ VGND VGND VPWR VPWR _12565_ sky130_fd_sc_hd__mux2_1
XFILLER_225_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25563_ _11063_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__clkbuf_1
X_22775_ _09410_ _09413_ _07369_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27302_ _12012_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24514_ _10476_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28282_ registers\[2\]\[20\] _10346_ _12528_ VGND VGND VPWR VPWR _12529_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21726_ registers\[36\]\[30\] registers\[37\]\[30\] registers\[38\]\[30\] registers\[39\]\[30\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__mux4_1
XFILLER_227_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25494_ _11027_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27233_ _11805_ registers\[37\]\[36\] _11969_ VGND VGND VPWR VPWR _11976_ sky130_fd_sc_hd__mux2_1
X_24445_ _10439_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__buf_4
XFILLER_8_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21657_ registers\[56\]\[28\] registers\[57\]\[28\] registers\[58\]\[28\] registers\[59\]\[28\]
+ _08194_ _08327_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__mux4_1
XFILLER_205_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_84_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_84_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20608_ registers\[36\]\[0\] registers\[37\]\[0\] registers\[38\]\[0\] registers\[39\]\[0\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__mux4_1
X_27164_ _11736_ registers\[37\]\[3\] _11936_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24376_ net37 VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21588_ registers\[60\]\[26\] registers\[61\]\[26\] registers\[62\]\[26\] registers\[63\]\[26\]
+ _08198_ _07992_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__mux4_1
X_26115_ _11300_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__buf_4
X_23327_ net53 VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__buf_4
X_20539_ registers\[28\]\[62\] registers\[29\]\[62\] registers\[30\]\[62\] registers\[31\]\[62\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__mux4_1
XFILLER_193_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27095_ _11903_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26046_ _10766_ registers\[45\]\[17\] _11312_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23258_ _09767_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22209_ registers\[24\]\[43\] registers\[25\]\[43\] registers\[26\]\[43\] registers\[27\]\[43\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__mux4_1
XTAP_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23189_ registers\[9\]\[12\] _09683_ _09722_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__mux2_1
XTAP_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1405 _00177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1416 _00181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1427 _04646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29805_ registers\[18\]\[7\] _12949_ _13353_ VGND VGND VPWR VPWR _13361_ sky130_fd_sc_hd__mux2_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1438 _05059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1449 _05073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27997_ _11757_ registers\[31\]\[13\] _12375_ VGND VGND VPWR VPWR _12379_ sky130_fd_sc_hd__mux2_1
XTAP_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17750_ _04294_ _04528_ _04529_ _04299_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__a22o_1
X_29736_ _13324_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__clkbuf_1
X_26948_ _11813_ registers\[3\]\[40\] _11814_ VGND VGND VPWR VPWR _11815_ sky130_fd_sc_hd__mux2_1
XTAP_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ _15193_ _15196_ _14926_ VGND VGND VPWR VPWR _15197_ sky130_fd_sc_hd__o21ba_1
XTAP_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29667_ _13288_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__clkbuf_1
X_17681_ _04459_ _04462_ _04301_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__o21ba_1
X_26879_ _11767_ registers\[3\]\[18\] _11751_ VGND VGND VPWR VPWR _11768_ sky130_fd_sc_hd__mux2_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19420_ registers\[40\]\[30\] registers\[41\]\[30\] registers\[42\]\[30\] registers\[43\]\[30\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__mux4_1
X_28618_ _12705_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16632_ registers\[56\]\[16\] registers\[57\]\[16\] registers\[58\]\[16\] registers\[59\]\[16\]
+ _15066_ _14856_ VGND VGND VPWR VPWR _15130_ sky130_fd_sc_hd__mux4_1
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29598_ registers\[20\]\[37\] _13012_ _13244_ VGND VGND VPWR VPWR _13252_ sky130_fd_sc_hd__mux2_1
X_19351_ registers\[44\]\[28\] registers\[45\]\[28\] registers\[46\]\[28\] registers\[47\]\[28\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__mux4_1
X_28549_ _11769_ registers\[27\]\[19\] _12659_ VGND VGND VPWR VPWR _12669_ sky130_fd_sc_hd__mux2_1
X_16563_ registers\[36\]\[14\] registers\[37\]\[14\] registers\[38\]\[14\] registers\[39\]\[14\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _15063_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18302_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__buf_12
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31560_ _14284_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16494_ _14567_ VGND VGND VPWR VPWR _14996_ sky130_fd_sc_hd__clkbuf_4
X_19282_ registers\[36\]\[26\] registers\[37\]\[26\] registers\[38\]\[26\] registers\[39\]\[26\]
+ _05713_ _05714_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__mux4_1
XFILLER_128_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18233_ registers\[4\]\[62\] registers\[5\]\[62\] registers\[6\]\[62\] registers\[7\]\[62\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux4_1
XFILLER_15_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30511_ _09702_ registers\[13\]\[21\] _13731_ VGND VGND VPWR VPWR _13733_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31491_ _09771_ registers\[6\]\[38\] _14239_ VGND VGND VPWR VPWR _14248_ sky130_fd_sc_hd__mux2_1
XFILLER_31_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_75_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30442_ _13696_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33230_ clknet_leaf_74_CLK _01344_ VGND VGND VPWR VPWR registers\[48\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18164_ _14587_ _04929_ _04930_ _14597_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__a22o_1
XFILLER_156_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17115_ registers\[20\]\[29\] registers\[21\]\[29\] registers\[22\]\[29\] registers\[23\]\[29\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15600_ sky130_fd_sc_hd__mux4_1
X_18095_ registers\[40\]\[58\] registers\[41\]\[58\] registers\[42\]\[58\] registers\[43\]\[58\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__mux4_1
X_33161_ clknet_leaf_209_CLK _01275_ VGND VGND VPWR VPWR registers\[50\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30373_ _13637_ VGND VGND VPWR VPWR _13660_ sky130_fd_sc_hd__buf_4
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32112_ clknet_leaf_468_CLK _00027_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dfxtp_1
X_17046_ _15511_ _15518_ _15525_ _15532_ VGND VGND VPWR VPWR _15533_ sky130_fd_sc_hd__or4_4
X_33092_ clknet_leaf_258_CLK _01206_ VGND VGND VPWR VPWR registers\[51\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32043_ clknet_leaf_422_CLK _00221_ VGND VGND VPWR VPWR registers\[62\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _05540_ _05740_ _05741_ _05545_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__a22o_1
XFILLER_225_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35802_ clknet_leaf_14_CLK _03916_ VGND VGND VPWR VPWR registers\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _04540_ _04720_ _04721_ _04546_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__a22o_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33994_ clknet_leaf_159_CLK _02108_ VGND VGND VPWR VPWR registers\[37\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35733_ clknet_leaf_104_CLK _03847_ VGND VGND VPWR VPWR registers\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_32945_ clknet_leaf_367_CLK _01059_ VGND VGND VPWR VPWR registers\[53\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17879_ registers\[48\]\[51\] registers\[49\]\[51\] registers\[50\]\[51\] registers\[51\]\[51\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__mux4_1
XFILLER_61_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_26__f_CLK clknet_5_13_0_CLK VGND VGND VPWR VPWR clknet_6_26__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19618_ registers\[12\]\[35\] registers\[13\]\[35\] registers\[14\]\[35\] registers\[15\]\[35\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__mux4_1
X_35664_ clknet_leaf_135_CLK _03778_ VGND VGND VPWR VPWR registers\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20890_ registers\[0\]\[6\] registers\[1\]\[6\] registers\[2\]\[6\] registers\[3\]\[6\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__mux4_1
X_32876_ clknet_leaf_373_CLK _00990_ VGND VGND VPWR VPWR registers\[54\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_34615_ clknet_leaf_311_CLK _02729_ VGND VGND VPWR VPWR registers\[27\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31827_ _09668_ registers\[49\]\[5\] _14419_ VGND VGND VPWR VPWR _14425_ sky130_fd_sc_hd__mux2_1
X_19549_ _06031_ _06277_ _06278_ _06034_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__a22o_1
X_35595_ clknet_leaf_150_CLK _03709_ VGND VGND VPWR VPWR registers\[12\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22560_ _08958_ _09204_ _09205_ _08961_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__a22o_1
X_34546_ clknet_leaf_386_CLK _02660_ VGND VGND VPWR VPWR registers\[28\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31758_ _14388_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21511_ _08186_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
X_30709_ registers\[12\]\[51\] _13042_ _13835_ VGND VGND VPWR VPWR _13837_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22491_ _09135_ _09138_ _09102_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34477_ clknet_leaf_388_CLK _02591_ VGND VGND VPWR VPWR registers\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_31689_ _14352_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_66_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_66_CLK sky130_fd_sc_hd__clkbuf_16
X_24230_ _09634_ registers\[58\]\[57\] _10288_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__mux2_1
X_36216_ clknet_leaf_115_CLK _00100_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33428_ clknet_leaf_125_CLK _01542_ VGND VGND VPWR VPWR registers\[45\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_21442_ _07312_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36147_ clknet_leaf_364_CLK _04261_ VGND VGND VPWR VPWR registers\[49\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_24161_ _09565_ registers\[58\]\[24\] _10255_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__mux2_1
X_33359_ clknet_leaf_130_CLK _01473_ VGND VGND VPWR VPWR registers\[46\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_839 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21373_ registers\[36\]\[20\] registers\[37\]\[20\] registers\[38\]\[20\] registers\[39\]\[20\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__mux4_1
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23112_ registers\[39\]\[8\] _09674_ _09658_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20324_ _06722_ _07030_ _07031_ _06725_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__a22o_1
X_24092_ _09632_ registers\[5\]\[56\] _10216_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__mux2_1
XFILLER_190_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36078_ clknet_leaf_371_CLK _04192_ VGND VGND VPWR VPWR registers\[59\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23043_ _09625_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
X_35029_ clknet_leaf_104_CLK _03143_ VGND VGND VPWR VPWR registers\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_27920_ _12338_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__clkbuf_1
X_20255_ _06717_ _06963_ _06964_ _06720_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__a22o_1
XFILLER_235_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27851_ registers\[32\]\[8\] _10321_ _12293_ VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__mux2_1
X_20186_ registers\[0\]\[51\] registers\[1\]\[51\] registers\[2\]\[51\] registers\[3\]\[51\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__mux4_1
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26802_ _11718_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__clkbuf_1
XTAP_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24994_ _10732_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__clkbuf_1
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27782_ _12265_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__clkbuf_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29521_ registers\[20\]\[0\] _12931_ _13211_ VGND VGND VPWR VPWR _13212_ sky130_fd_sc_hd__mux2_1
XFILLER_170_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23945_ _10145_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26733_ _11682_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26664_ _11645_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29452_ _13175_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_803 _08973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23876_ _09552_ registers\[60\]\[18\] _10100_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__mux2_1
XANTENNA_814 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_825 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_836 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25615_ _11092_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
X_28403_ _12592_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22827_ _07385_ _09462_ _09463_ _07395_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__a22o_1
XFILLER_189_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_847 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29383_ _13138_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26595_ _11609_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_858 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_869 _09393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28334_ registers\[2\]\[45\] _10399_ _12550_ VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__mux2_1
XFILLER_129_1362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25546_ _11054_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22758_ registers\[44\]\[60\] registers\[45\]\[60\] registers\[46\]\[60\] registers\[47\]\[60\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__mux4_1
XFILLER_73_1136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21709_ _08272_ _08377_ _08378_ _08275_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__a22o_1
X_28265_ registers\[2\]\[12\] _10330_ _12517_ VGND VGND VPWR VPWR _12520_ sky130_fd_sc_hd__mux2_1
X_25477_ _11018_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22689_ registers\[28\]\[57\] registers\[29\]\[57\] registers\[30\]\[57\] registers\[31\]\[57\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_57_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_57_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24428_ net55 VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__buf_4
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27216_ _11788_ registers\[37\]\[28\] _11958_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__mux2_1
X_28196_ _12483_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27147_ _11930_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24359_ _10381_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27078_ _11894_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__clkbuf_1
X_26029_ _10749_ registers\[45\]\[9\] _11301_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__mux2_1
X_18920_ registers\[20\]\[15\] registers\[21\]\[15\] registers\[22\]\[15\] registers\[23\]\[15\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__mux4_1
XTAP_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1202 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1213 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18851_ registers\[16\]\[13\] registers\[17\]\[13\] registers\[18\]\[13\] registers\[19\]\[13\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__mux4_1
XTAP_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1224 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1235 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1246 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17802_ _04576_ _04579_ _15955_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1257 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1268 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18782_ _05496_ _05532_ _05533_ _05499_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__a22o_1
XFILLER_95_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1279 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15994_ net67 net68 VGND VGND VPWR VPWR _14508_ sky130_fd_sc_hd__and2_1
XTAP_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _15884_ _04511_ _04512_ _15890_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__a22o_1
X_29719_ registers\[1\]\[30\] _12997_ _13315_ VGND VGND VPWR VPWR _13316_ sky130_fd_sc_hd__mux2_1
XFILLER_236_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30991_ registers\[10\]\[57\] _13054_ _13977_ VGND VGND VPWR VPWR _13985_ sky130_fd_sc_hd__mux2_1
XTAP_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32730_ clknet_leaf_68_CLK _00844_ VGND VGND VPWR VPWR registers\[56\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17664_ _15892_ _04444_ _04445_ _15896_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a22o_1
XFILLER_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19403_ _06133_ _06136_ _05826_ _05827_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__o211a_1
X_16615_ _15110_ _15113_ _14945_ VGND VGND VPWR VPWR _15114_ sky130_fd_sc_hd__o21ba_1
X_32661_ clknet_leaf_69_CLK _00775_ VGND VGND VPWR VPWR registers\[57\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17595_ _15884_ _04377_ _04378_ _15890_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a22o_1
XFILLER_189_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34400_ clknet_leaf_490_CLK _02514_ VGND VGND VPWR VPWR registers\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19334_ _06031_ _06068_ _06069_ _06034_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__a22o_1
X_31612_ registers\[63\]\[31\] net25 _14310_ VGND VGND VPWR VPWR _14312_ sky130_fd_sc_hd__mux2_1
X_16546_ registers\[12\]\[13\] registers\[13\]\[13\] registers\[14\]\[13\] registers\[15\]\[13\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15047_ sky130_fd_sc_hd__mux4_1
X_35380_ clknet_leaf_416_CLK _03494_ VGND VGND VPWR VPWR registers\[15\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32592_ clknet_leaf_75_CLK _00706_ VGND VGND VPWR VPWR registers\[58\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34331_ clknet_leaf_1_CLK _02445_ VGND VGND VPWR VPWR registers\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_31543_ _09825_ registers\[6\]\[63\] _14205_ VGND VGND VPWR VPWR _14275_ sky130_fd_sc_hd__mux2_1
X_19265_ registers\[12\]\[25\] registers\[13\]\[25\] registers\[14\]\[25\] registers\[15\]\[25\]
+ _05937_ _05938_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__mux4_1
X_16477_ registers\[4\]\[11\] registers\[5\]\[11\] registers\[6\]\[11\] registers\[7\]\[11\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _14980_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_48_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_48_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18216_ registers\[32\]\[62\] registers\[33\]\[62\] registers\[34\]\[62\] registers\[35\]\[62\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__mux4_1
X_34262_ clknet_leaf_124_CLK _02376_ VGND VGND VPWR VPWR registers\[32\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_19196_ _05688_ _05934_ _05935_ _05691_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a22o_1
XFILLER_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31474_ _14205_ VGND VGND VPWR VPWR _14239_ sky130_fd_sc_hd__buf_6
XFILLER_191_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36001_ clknet_leaf_444_CLK _04115_ VGND VGND VPWR VPWR registers\[63\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33213_ clknet_leaf_305_CLK _01327_ VGND VGND VPWR VPWR registers\[4\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_18147_ registers\[16\]\[59\] registers\[17\]\[59\] registers\[18\]\[59\] registers\[19\]\[59\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__mux4_1
X_30425_ _13687_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__clkbuf_1
X_34193_ clknet_leaf_129_CLK _02307_ VGND VGND VPWR VPWR registers\[33\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33144_ clknet_leaf_333_CLK _01258_ VGND VGND VPWR VPWR registers\[50\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_18078_ _04844_ _04847_ _04619_ _04620_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__o211a_1
X_30356_ _13651_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17029_ registers\[52\]\[27\] registers\[53\]\[27\] registers\[54\]\[27\] registers\[55\]\[27\]
+ _15477_ _15478_ VGND VGND VPWR VPWR _15516_ sky130_fd_sc_hd__mux4_1
XFILLER_217_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30287_ _13614_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__clkbuf_1
X_33075_ clknet_leaf_358_CLK _01189_ VGND VGND VPWR VPWR registers\[51\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_20040_ _06717_ _06754_ _06755_ _06720_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__a22o_1
XFILLER_193_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32026_ clknet_leaf_66_CLK _00204_ VGND VGND VPWR VPWR registers\[62\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1780 _12718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1791 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33977_ clknet_leaf_281_CLK _02091_ VGND VGND VPWR VPWR registers\[37\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21991_ _08649_ _08652_ _08416_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35716_ clknet_leaf_225_CLK _03830_ VGND VGND VPWR VPWR registers\[10\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23730_ _09542_ registers\[29\]\[13\] _10028_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__mux2_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ registers\[40\]\[8\] registers\[41\]\[8\] registers\[42\]\[8\] registers\[43\]\[8\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__mux4_1
XFILLER_54_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32928_ clknet_leaf_45_CLK _01042_ VGND VGND VPWR VPWR registers\[53\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35647_ clknet_leaf_296_CLK _03761_ VGND VGND VPWR VPWR registers\[11\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_23661_ registers\[61\]\[46\] _09788_ _09987_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__mux2_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20873_ registers\[32\]\[6\] registers\[33\]\[6\] registers\[34\]\[6\] registers\[35\]\[6\]
+ _07304_ _07306_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__mux4_1
X_32859_ clknet_leaf_54_CLK _00973_ VGND VGND VPWR VPWR registers\[54\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_25400_ _10804_ registers\[50\]\[35\] _10970_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__mux2_1
X_22612_ registers\[56\]\[55\] registers\[57\]\[55\] registers\[58\]\[55\] registers\[59\]\[55\]
+ _09223_ _09013_ VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__mux4_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26380_ _11495_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35578_ clknet_leaf_302_CLK _03692_ VGND VGND VPWR VPWR registers\[12\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_23592_ registers\[61\]\[13\] _09685_ _09954_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__mux2_1
XFILLER_74_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25331_ _10735_ registers\[50\]\[2\] _10937_ VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__mux2_1
XFILLER_224_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22543_ registers\[36\]\[53\] registers\[37\]\[53\] registers\[38\]\[53\] registers\[39\]\[53\]
+ _08978_ _08979_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__mux4_1
XFILLER_210_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34529_ clknet_leaf_488_CLK _02643_ VGND VGND VPWR VPWR registers\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_39_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_39_CLK sky130_fd_sc_hd__clkbuf_16
X_28050_ _12406_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25262_ _10802_ registers\[51\]\[34\] _10898_ VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__mux2_1
X_22474_ registers\[44\]\[51\] registers\[45\]\[51\] registers\[46\]\[51\] registers\[47\]\[51\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__mux4_1
X_27001_ _11850_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_1
X_24213_ _09617_ registers\[58\]\[49\] _10277_ VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__mux2_1
X_21425_ _08099_ _08102_ _08062_ _08063_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__o211a_1
X_25193_ _10733_ registers\[51\]\[1\] _10865_ VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__mux2_1
XFILLER_198_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24144_ _09548_ registers\[58\]\[16\] _10244_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__mux2_1
XFILLER_136_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21356_ _07929_ _08034_ _08035_ _07932_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__a22o_1
XFILLER_136_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20307_ _06912_ _07013_ _07014_ _06917_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__a22o_1
XFILLER_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24075_ _09615_ registers\[5\]\[48\] _10205_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__mux2_1
XFILLER_151_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28952_ registers\[24\]\[18\] _10342_ _12872_ VGND VGND VPWR VPWR _12881_ sky130_fd_sc_hd__mux2_1
X_21287_ registers\[16\]\[17\] registers\[17\]\[17\] registers\[18\]\[17\] registers\[19\]\[17\]
+ _07936_ _07937_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__mux4_1
X_23026_ _09613_ registers\[62\]\[47\] _09599_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__mux2_1
XFILLER_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27903_ _12329_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20238_ _06948_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__buf_4
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28883_ _12844_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27834_ _12292_ VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__buf_6
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20169_ _06848_ _06857_ _06867_ _06881_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__or4_2
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27765_ registers\[33\]\[31\] _10370_ _12255_ VGND VGND VPWR VPWR _12257_ sky130_fd_sc_hd__mux2_1
X_24977_ _09636_ registers\[53\]\[58\] _10713_ VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__mux2_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29504_ _13202_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__clkbuf_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26716_ _11673_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ _10136_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_218_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27696_ registers\[34\]\[63\] _10436_ _12150_ VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__mux2_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_600 _05088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_611 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_622 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29435_ _13166_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__clkbuf_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26647_ _11636_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_633 _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23859_ _10088_ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__clkbuf_8
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_644 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_655 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_666 _05396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16400_ _14796_ _14903_ _14904_ _14799_ VGND VGND VPWR VPWR _14905_ sky130_fd_sc_hd__a22o_1
XFILLER_60_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29366_ _09808_ registers\[22\]\[55\] _13124_ VGND VGND VPWR VPWR _13130_ sky130_fd_sc_hd__mux2_1
XANTENNA_677 _05853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17380_ _15541_ _15855_ _15856_ _15547_ VGND VGND VPWR VPWR _15857_ sky130_fd_sc_hd__a22o_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_688 _06300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26578_ _11600_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_699 _07275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16331_ _14801_ _14836_ _14837_ _14804_ VGND VGND VPWR VPWR _14838_ sky130_fd_sc_hd__a22o_1
X_28317_ registers\[2\]\[37\] _10382_ _12539_ VGND VGND VPWR VPWR _12547_ sky130_fd_sc_hd__mux2_1
X_25529_ registers\[4\]\[30\] _10367_ _11045_ VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__mux2_1
X_29297_ _09717_ registers\[22\]\[22\] _13091_ VGND VGND VPWR VPWR _13094_ sky130_fd_sc_hd__mux2_1
XFILLER_13_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16262_ _14767_ _14770_ _14585_ VGND VGND VPWR VPWR _14771_ sky130_fd_sc_hd__o21ba_1
X_19050_ _05790_ _05793_ _05483_ _05484_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__o211a_1
XFILLER_200_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28248_ registers\[2\]\[4\] _10313_ _12506_ VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__mux2_1
XFILLER_139_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18001_ _04637_ _04772_ _04773_ _04642_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__a22o_1
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16193_ registers\[12\]\[3\] registers\[13\]\[3\] registers\[14\]\[3\] registers\[15\]\[3\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14704_ sky130_fd_sc_hd__mux4_1
XFILLER_12_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28179_ _12474_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30210_ registers\[15\]\[7\] _12949_ _13566_ VGND VGND VPWR VPWR _13574_ sky130_fd_sc_hd__mux2_1
XFILLER_138_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31190_ registers\[8\]\[23\] net16 _14086_ VGND VGND VPWR VPWR _14090_ sky130_fd_sc_hd__mux2_1
XFILLER_86_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30141_ _13537_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19952_ registers\[40\]\[45\] registers\[41\]\[45\] registers\[42\]\[45\] registers\[43\]\[45\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__mux4_1
XFILLER_218_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18903_ registers\[60\]\[15\] registers\[61\]\[15\] registers\[62\]\[15\] registers\[63\]\[15\]
+ _05619_ _05413_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__mux4_1
X_30072_ _13501_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__clkbuf_1
X_19883_ _06598_ _06603_ _06537_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1010 _11935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1021 _12505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1032 _12934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33900_ clknet_leaf_325_CLK _02014_ VGND VGND VPWR VPWR registers\[38\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1043 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18834_ registers\[56\]\[13\] registers\[57\]\[13\] registers\[58\]\[13\] registers\[59\]\[13\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__mux4_1
XTAP_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34880_ clknet_leaf_203_CLK _02994_ VGND VGND VPWR VPWR registers\[23\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1054 _13494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1065 _14063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1076 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1087 _14502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33831_ clknet_leaf_457_CLK _01945_ VGND VGND VPWR VPWR registers\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1098 _14527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18765_ _05513_ _05516_ _05475_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__o21ba_1
X_15977_ _14490_ VGND VGND VPWR VPWR _14491_ sky130_fd_sc_hd__clkbuf_4
XTAP_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17716_ registers\[28\]\[46\] registers\[29\]\[46\] registers\[30\]\[46\] registers\[31\]\[46\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__mux4_1
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33762_ clknet_leaf_55_CLK _01876_ VGND VGND VPWR VPWR registers\[40\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_30974_ registers\[10\]\[49\] _13037_ _13966_ VGND VGND VPWR VPWR _13976_ sky130_fd_sc_hd__mux2_1
X_18696_ _05412_ _05448_ _05449_ _05416_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__a22o_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35501_ clknet_leaf_392_CLK _03615_ VGND VGND VPWR VPWR registers\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_32713_ clknet_leaf_209_CLK _00827_ VGND VGND VPWR VPWR registers\[57\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_17647_ registers\[20\]\[44\] registers\[21\]\[44\] registers\[22\]\[44\] registers\[23\]\[44\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__mux4_1
XFILLER_64_987 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_224_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33693_ clknet_leaf_28_CLK _01807_ VGND VGND VPWR VPWR registers\[41\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35432_ clknet_leaf_399_CLK _03546_ VGND VGND VPWR VPWR registers\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_32644_ clknet_leaf_264_CLK _00758_ VGND VGND VPWR VPWR registers\[58\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_17578_ _14576_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__buf_6
XFILLER_56_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19317_ registers\[32\]\[27\] registers\[33\]\[27\] registers\[34\]\[27\] registers\[35\]\[27\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__mux4_1
X_35363_ clknet_leaf_469_CLK _03477_ VGND VGND VPWR VPWR registers\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_16529_ _14991_ _15028_ _15029_ _14996_ VGND VGND VPWR VPWR _15030_ sky130_fd_sc_hd__a22o_1
X_32575_ clknet_leaf_295_CLK _00689_ VGND VGND VPWR VPWR registers\[5\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34314_ clknet_leaf_156_CLK _02428_ VGND VGND VPWR VPWR registers\[32\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_31526_ _14266_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__clkbuf_1
X_19248_ _05883_ _05984_ _05985_ _05888_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__a22o_1
XFILLER_177_878 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35294_ clknet_leaf_3_CLK _03408_ VGND VGND VPWR VPWR registers\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34245_ clknet_leaf_245_CLK _02359_ VGND VGND VPWR VPWR registers\[33\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_31457_ _14230_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__clkbuf_1
X_19179_ _05919_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__clkbuf_1
X_21210_ registers\[0\]\[15\] registers\[1\]\[15\] registers\[2\]\[15\] registers\[3\]\[15\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__mux4_1
X_30408_ _13678_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__clkbuf_1
X_34176_ clknet_leaf_258_CLK _02290_ VGND VGND VPWR VPWR registers\[34\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_22190_ registers\[36\]\[43\] registers\[37\]\[43\] registers\[38\]\[43\] registers\[39\]\[43\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__mux4_1
X_31388_ registers\[7\]\[53\] net49 _14190_ VGND VGND VPWR VPWR _14194_ sky130_fd_sc_hd__mux2_1
XFILLER_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_5_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_5_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21141_ registers\[8\]\[13\] registers\[9\]\[13\] registers\[10\]\[13\] registers\[11\]\[13\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__mux4_1
X_33127_ clknet_leaf_434_CLK _01241_ VGND VGND VPWR VPWR registers\[50\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_30339_ _13642_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21072_ _07756_ _07759_ _07719_ _07720_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__o211a_1
X_33058_ clknet_leaf_46_CLK _01172_ VGND VGND VPWR VPWR registers\[51\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20023_ registers\[32\]\[47\] registers\[33\]\[47\] registers\[34\]\[47\] registers\[35\]\[47\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__mux4_1
X_32009_ clknet_leaf_29_CLK _00182_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24900_ _09559_ registers\[53\]\[21\] _10680_ VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__mux2_1
X_25880_ _10735_ registers\[46\]\[2\] _11230_ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__mux2_1
XFILLER_140_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24831_ _10645_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27550_ _12142_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__clkbuf_1
X_24762_ _10586_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__buf_4
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21974_ _07358_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__clkbuf_4
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23713_ _09525_ registers\[29\]\[5\] _10017_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__mux2_1
X_26501_ _11559_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__clkbuf_1
X_20925_ _07613_ _07616_ _07339_ _07341_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__o211a_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27481_ _12106_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__clkbuf_1
X_24693_ _09624_ registers\[55\]\[52\] _10569_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__mux2_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29220_ registers\[23\]\[54\] _13048_ _13040_ VGND VGND VPWR VPWR _13049_ sky130_fd_sc_hd__mux2_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26432_ _10747_ registers\[42\]\[8\] _11514_ VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__mux2_1
XFILLER_230_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_199_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23644_ registers\[61\]\[38\] _09771_ _09976_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__mux2_1
X_20856_ registers\[8\]\[5\] registers\[9\]\[5\] registers\[10\]\[5\] registers\[11\]\[5\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__mux4_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29151_ net26 VGND VGND VPWR VPWR _13002_ sky130_fd_sc_hd__clkbuf_4
X_26363_ _11486_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23575_ registers\[61\]\[5\] _09668_ _09943_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__mux2_1
X_20787_ _07479_ _07482_ _07339_ _07341_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__o211a_1
X_28102_ _12433_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__clkbuf_1
X_25314_ _10854_ registers\[51\]\[59\] _10920_ VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__mux2_1
X_22526_ _08958_ _09171_ _09172_ _08961_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__a22o_1
X_26294_ _11450_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29082_ net2 VGND VGND VPWR VPWR _12955_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28033_ _11792_ registers\[31\]\[30\] _12397_ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__mux2_1
X_25245_ _10785_ registers\[51\]\[26\] _10887_ VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__mux2_1
X_22457_ registers\[16\]\[50\] registers\[17\]\[50\] registers\[18\]\[50\] registers\[19\]\[50\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__mux4_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21408_ _07398_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__buf_2
X_25176_ _10855_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22388_ registers\[28\]\[48\] registers\[29\]\[48\] registers\[30\]\[48\] registers\[31\]\[48\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__mux4_1
X_24127_ _09531_ registers\[58\]\[8\] _10233_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__mux2_1
XFILLER_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21339_ _07776_ _08015_ _08018_ _07781_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__a22o_1
XFILLER_124_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29984_ registers\[17\]\[28\] _12993_ _13446_ VGND VGND VPWR VPWR _13455_ sky130_fd_sc_hd__mux2_1
XFILLER_151_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24058_ _10160_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__buf_4
X_28935_ net282 VGND VGND VPWR VPWR _12872_ sky130_fd_sc_hd__buf_4
XFILLER_137_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23009_ _09602_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28866_ _11816_ registers\[25\]\[41\] _12834_ VGND VGND VPWR VPWR _12836_ sky130_fd_sc_hd__mux2_1
X_16880_ registers\[40\]\[23\] registers\[41\]\[23\] registers\[42\]\[23\] registers\[43\]\[23\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15371_ sky130_fd_sc_hd__mux4_1
XFILLER_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27817_ registers\[33\]\[56\] _10422_ _12277_ VGND VGND VPWR VPWR _12284_ sky130_fd_sc_hd__mux2_1
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28797_ _12799_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__clkbuf_1
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18550_ registers\[60\]\[5\] registers\[61\]\[5\] registers\[62\]\[5\] registers\[63\]\[5\]
+ _05276_ _05093_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__mux4_1
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27748_ registers\[33\]\[23\] _10353_ _12244_ VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__mux2_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17501_ _15970_ _15973_ _15974_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__o21ba_1
XFILLER_205_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ registers\[56\]\[3\] registers\[57\]\[3\] registers\[58\]\[3\] registers\[59\]\[3\]
+ _05079_ _05081_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__mux4_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27679_ _12211_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_430 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_441 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29418_ _13157_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17432_ registers\[24\]\[38\] registers\[25\]\[38\] registers\[26\]\[38\] registers\[27\]\[38\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15908_ sky130_fd_sc_hd__mux4_1
XANTENNA_452 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_463 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_474 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30690_ registers\[12\]\[42\] _13023_ _13824_ VGND VGND VPWR VPWR _13827_ sky130_fd_sc_hd__mux2_1
XFILLER_198_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_496 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29349_ _09791_ registers\[22\]\[47\] _13113_ VGND VGND VPWR VPWR _13121_ sky130_fd_sc_hd__mux2_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17363_ registers\[28\]\[36\] registers\[29\]\[36\] registers\[30\]\[36\] registers\[31\]\[36\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15841_ sky130_fd_sc_hd__mux4_1
XFILLER_186_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19102_ registers\[28\]\[20\] registers\[29\]\[20\] registers\[30\]\[20\] registers\[31\]\[20\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__mux4_1
XFILLER_105_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16314_ _14571_ VGND VGND VPWR VPWR _14821_ sky130_fd_sc_hd__buf_6
XFILLER_242_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32360_ clknet_leaf_436_CLK _00474_ VGND VGND VPWR VPWR registers\[61\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17294_ registers\[20\]\[34\] registers\[21\]\[34\] registers\[22\]\[34\] registers\[23\]\[34\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15774_ sky130_fd_sc_hd__mux4_1
XFILLER_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19033_ _05746_ _05761_ _05770_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__or4_1
X_31311_ _14153_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16245_ _14655_ _14752_ _14753_ _14658_ VGND VGND VPWR VPWR _14754_ sky130_fd_sc_hd__a22o_1
X_32291_ clknet_leaf_474_CLK _00405_ VGND VGND VPWR VPWR registers\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34030_ clknet_leaf_359_CLK _02144_ VGND VGND VPWR VPWR registers\[36\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_31242_ registers\[8\]\[48\] net43 _14108_ VGND VGND VPWR VPWR _14117_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16176_ _14648_ _14685_ _14686_ _14653_ VGND VGND VPWR VPWR _14687_ sky130_fd_sc_hd__a22o_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput106 net106 VGND VGND VPWR VPWR D1[24] sky130_fd_sc_hd__buf_2
XFILLER_182_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput117 net117 VGND VGND VPWR VPWR D1[34] sky130_fd_sc_hd__buf_2
Xoutput128 net128 VGND VGND VPWR VPWR D1[44] sky130_fd_sc_hd__buf_2
XFILLER_142_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput139 net139 VGND VGND VPWR VPWR D1[54] sky130_fd_sc_hd__buf_2
X_31173_ registers\[8\]\[15\] net7 _14075_ VGND VGND VPWR VPWR _14081_ sky130_fd_sc_hd__mux2_1
XFILLER_181_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19935_ registers\[0\]\[44\] registers\[1\]\[44\] registers\[2\]\[44\] registers\[3\]\[44\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__mux4_1
X_30124_ registers\[16\]\[30\] _12997_ _13528_ VGND VGND VPWR VPWR _13529_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35981_ clknet_leaf_145_CLK _04095_ VGND VGND VPWR VPWR registers\[6\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30055_ registers\[17\]\[62\] _13064_ _13423_ VGND VGND VPWR VPWR _13492_ sky130_fd_sc_hd__mux2_1
X_34932_ clknet_leaf_414_CLK _03046_ VGND VGND VPWR VPWR registers\[22\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_19866_ _06441_ _06585_ _06586_ _06445_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__a22o_1
XFILLER_214_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_233_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18817_ registers\[16\]\[12\] registers\[17\]\[12\] registers\[18\]\[12\] registers\[19\]\[12\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__mux4_1
X_34863_ clknet_leaf_395_CLK _02977_ VGND VGND VPWR VPWR registers\[23\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19797_ registers\[12\]\[40\] registers\[13\]\[40\] registers\[14\]\[40\] registers\[15\]\[40\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__mux4_1
XFILLER_231_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33814_ clknet_leaf_88_CLK _01928_ VGND VGND VPWR VPWR registers\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_18748_ _05149_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34794_ clknet_leaf_451_CLK _02908_ VGND VGND VPWR VPWR registers\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33745_ clknet_leaf_130_CLK _01859_ VGND VGND VPWR VPWR registers\[40\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_18679_ _05430_ _05433_ _05163_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__o21ba_1
XFILLER_63_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30957_ _13967_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20710_ registers\[36\]\[1\] registers\[37\]\[1\] registers\[38\]\[1\] registers\[39\]\[1\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__mux4_1
XFILLER_149_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33676_ clknet_leaf_171_CLK _01790_ VGND VGND VPWR VPWR registers\[42\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_21690_ _07305_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__buf_4
XFILLER_180_1109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30888_ registers\[10\]\[8\] _12951_ _13922_ VGND VGND VPWR VPWR _13931_ sky130_fd_sc_hd__mux2_1
XFILLER_196_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35415_ clknet_leaf_82_CLK _03529_ VGND VGND VPWR VPWR registers\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_20641_ net76 VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__buf_12
X_32627_ clknet_leaf_363_CLK _00741_ VGND VGND VPWR VPWR registers\[58\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35346_ clknet_leaf_77_CLK _03460_ VGND VGND VPWR VPWR registers\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_23360_ _09833_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
X_20572_ _07268_ _07271_ _05162_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__o21ba_1
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32558_ clknet_leaf_376_CLK _00672_ VGND VGND VPWR VPWR registers\[5\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22311_ registers\[24\]\[46\] registers\[25\]\[46\] registers\[26\]\[46\] registers\[27\]\[46\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__mux4_1
XFILLER_178_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31509_ _14257_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35277_ clknet_leaf_148_CLK _03391_ VGND VGND VPWR VPWR registers\[17\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23291_ _09789_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32489_ clknet_leaf_407_CLK _00603_ VGND VGND VPWR VPWR registers\[60\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25030_ _10756_ registers\[52\]\[12\] _10752_ VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__mux2_1
X_22242_ _07349_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__clkbuf_8
XFILLER_178_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34228_ clknet_leaf_349_CLK _02342_ VGND VGND VPWR VPWR registers\[33\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22173_ _08615_ _08828_ _08829_ _08618_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__a22o_1
X_34159_ clknet_leaf_355_CLK _02273_ VGND VGND VPWR VPWR registers\[34\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21124_ _07805_ _07810_ _07744_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__o21ba_1
XFILLER_105_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26981_ net47 VGND VGND VPWR VPWR _11837_ sky130_fd_sc_hd__buf_4
XFILLER_120_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28720_ _11805_ registers\[26\]\[36\] _12752_ VGND VGND VPWR VPWR _12759_ sky130_fd_sc_hd__mux2_1
X_25932_ _10787_ registers\[46\]\[27\] _11252_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21055_ _07398_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__buf_2
XFILLER_232_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20006_ registers\[12\]\[46\] registers\[13\]\[46\] registers\[14\]\[46\] registers\[15\]\[46\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__mux4_1
XFILLER_219_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28651_ _11736_ registers\[26\]\[3\] _12719_ VGND VGND VPWR VPWR _12723_ sky130_fd_sc_hd__mux2_1
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25863_ _11223_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27602_ registers\[34\]\[18\] _10342_ _12162_ VGND VGND VPWR VPWR _12171_ sky130_fd_sc_hd__mux2_1
XFILLER_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24814_ _10636_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28582_ _12686_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__clkbuf_1
X_25794_ _11187_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ _11834_ registers\[35\]\[50\] _12133_ VGND VGND VPWR VPWR _12134_ sky130_fd_sc_hd__mux2_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24745_ _10600_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
X_21957_ _08614_ _08619_ _08416_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__o21ba_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_270_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_270_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _07571_ _07580_ _07591_ _07600_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__or4_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24676_ _09607_ registers\[55\]\[44\] _10558_ VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__mux2_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27464_ _12097_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__clkbuf_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21888_ _07347_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__buf_6
XFILLER_203_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29203_ net44 VGND VGND VPWR VPWR _13037_ sky130_fd_sc_hd__clkbuf_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26415_ _11513_ VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__buf_4
XFILLER_208_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23627_ _09942_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__buf_4
XFILLER_208_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20839_ _07533_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27395_ registers\[36\]\[49\] _10407_ _12051_ VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__mux2_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29134_ _12990_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__clkbuf_1
X_23558_ _09938_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26346_ _10796_ registers\[43\]\[31\] _11476_ VGND VGND VPWR VPWR _11478_ sky130_fd_sc_hd__mux2_1
XFILLER_11_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22509_ registers\[44\]\[52\] registers\[45\]\[52\] registers\[46\]\[52\] registers\[47\]\[52\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__mux4_1
XFILLER_155_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 DW[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_4
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26277_ _10862_ registers\[44\]\[63\] _11371_ VGND VGND VPWR VPWR _11441_ sky130_fd_sc_hd__mux2_1
X_29065_ registers\[23\]\[4\] _12943_ _12935_ VGND VGND VPWR VPWR _12944_ sky130_fd_sc_hd__mux2_1
X_23489_ _09902_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16030_ _14543_ VGND VGND VPWR VPWR _14544_ sky130_fd_sc_hd__buf_4
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28016_ _11776_ registers\[31\]\[22\] _12386_ VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25228_ _10768_ registers\[51\]\[18\] _10876_ VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__mux2_1
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25159_ net50 VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__buf_2
XFILLER_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17981_ _04540_ _04752_ _04753_ _04546_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__a22o_1
X_29967_ _13423_ VGND VGND VPWR VPWR _13446_ sky130_fd_sc_hd__buf_4
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19720_ _05065_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__clkbuf_4
X_28918_ _12863_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__clkbuf_1
X_16932_ registers\[4\]\[24\] registers\[5\]\[24\] registers\[6\]\[24\] registers\[7\]\[24\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15422_ sky130_fd_sc_hd__mux4_1
XFILLER_133_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29898_ registers\[18\]\[51\] _13042_ _13408_ VGND VGND VPWR VPWR _13410_ sky130_fd_sc_hd__mux2_1
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19651_ _06374_ _06375_ _06376_ _06377_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__a22o_1
X_16863_ registers\[0\]\[22\] registers\[1\]\[22\] registers\[2\]\[22\] registers\[3\]\[22\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15355_ sky130_fd_sc_hd__mux4_1
X_28849_ _11799_ registers\[25\]\[33\] _12823_ VGND VGND VPWR VPWR _12827_ sky130_fd_sc_hd__mux2_1
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18602_ registers\[16\]\[6\] registers\[17\]\[6\] registers\[18\]\[6\] registers\[19\]\[6\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__mux4_1
XFILLER_150_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19582_ registers\[0\]\[34\] registers\[1\]\[34\] registers\[2\]\[34\] registers\[3\]\[34\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux4_1
XFILLER_37_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31860_ _14442_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16794_ _14584_ VGND VGND VPWR VPWR _15288_ sky130_fd_sc_hd__buf_2
XFILLER_93_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_246_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18533_ _05137_ _05290_ _05291_ _05147_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__a22o_1
X_30811_ _13890_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_1242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31791_ registers\[59\]\[52\] net48 _14403_ VGND VGND VPWR VPWR _14406_ sky130_fd_sc_hd__mux2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_261_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_261_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_907 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33530_ clknet_leaf_279_CLK _01644_ VGND VGND VPWR VPWR registers\[44\]\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30742_ _13854_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__clkbuf_1
X_18464_ registers\[16\]\[2\] registers\[17\]\[2\] registers\[18\]\[2\] registers\[19\]\[2\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__mux4_1
XFILLER_34_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17415_ _15884_ _15886_ _15889_ _15890_ VGND VGND VPWR VPWR _15891_ sky130_fd_sc_hd__a22o_1
XANTENNA_293 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33461_ clknet_leaf_344_CLK _01575_ VGND VGND VPWR VPWR registers\[45\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_18395_ registers\[20\]\[0\] registers\[21\]\[0\] registers\[22\]\[0\] registers\[23\]\[0\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__mux4_1
X_30673_ registers\[12\]\[34\] _13006_ _13813_ VGND VGND VPWR VPWR _13818_ sky130_fd_sc_hd__mux2_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35200_ clknet_leaf_221_CLK _03314_ VGND VGND VPWR VPWR registers\[18\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32412_ clknet_leaf_0_CLK _00526_ VGND VGND VPWR VPWR registers\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_36180_ clknet_leaf_93_CLK _00124_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dfxtp_1
X_17346_ _15818_ _15823_ _15620_ _15621_ VGND VGND VPWR VPWR _15824_ sky130_fd_sc_hd__o211a_1
X_33392_ clknet_leaf_362_CLK _01506_ VGND VGND VPWR VPWR registers\[46\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35131_ clknet_leaf_301_CLK _03245_ VGND VGND VPWR VPWR registers\[1\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_32343_ clknet_leaf_61_CLK _00457_ VGND VGND VPWR VPWR registers\[61\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17277_ registers\[60\]\[34\] registers\[61\]\[34\] registers\[62\]\[34\] registers\[63\]\[34\]
+ _15756_ _15550_ VGND VGND VPWR VPWR _15757_ sky130_fd_sc_hd__mux4_1
XFILLER_228_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ _05754_ _05760_ _05483_ _05484_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__o211a_1
XFILLER_228_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16228_ _14734_ _14737_ _14585_ VGND VGND VPWR VPWR _14738_ sky130_fd_sc_hd__o21ba_1
X_35062_ clknet_leaf_304_CLK _03176_ VGND VGND VPWR VPWR registers\[20\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_32274_ clknet_leaf_101_CLK _00388_ VGND VGND VPWR VPWR registers\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34013_ clknet_leaf_26_CLK _02127_ VGND VGND VPWR VPWR registers\[36\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_31225_ _14063_ VGND VGND VPWR VPWR _14108_ sky130_fd_sc_hd__buf_4
XFILLER_114_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16159_ registers\[12\]\[2\] registers\[13\]\[2\] registers\[14\]\[2\] registers\[15\]\[2\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _14671_ sky130_fd_sc_hd__mux4_1
XFILLER_6_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31156_ registers\[8\]\[7\] net62 _14064_ VGND VGND VPWR VPWR _14072_ sky130_fd_sc_hd__mux2_1
XFILLER_142_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30107_ registers\[16\]\[22\] _12981_ _13517_ VGND VGND VPWR VPWR _13520_ sky130_fd_sc_hd__mux2_1
X_19918_ registers\[40\]\[44\] registers\[41\]\[44\] registers\[42\]\[44\] registers\[43\]\[44\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__mux4_1
XFILLER_155_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35964_ clknet_leaf_305_CLK _04078_ VGND VGND VPWR VPWR registers\[6\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31087_ _14035_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30038_ _13483_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__clkbuf_1
X_19849_ _05042_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__buf_4
XFILLER_29_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34915_ clknet_leaf_473_CLK _03029_ VGND VGND VPWR VPWR registers\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35895_ clknet_leaf_313_CLK _04009_ VGND VGND VPWR VPWR registers\[7\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22860_ registers\[0\]\[63\] registers\[1\]\[63\] registers\[2\]\[63\] registers\[3\]\[63\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__mux4_1
XFILLER_216_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34846_ clknet_leaf_491_CLK _02960_ VGND VGND VPWR VPWR registers\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21811_ registers\[60\]\[32\] registers\[61\]\[32\] registers\[62\]\[32\] registers\[63\]\[32\]
+ _08198_ _08335_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__mux4_1
XFILLER_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22791_ _09425_ _09428_ _07309_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__o21ba_1
X_34777_ clknet_leaf_20_CLK _02891_ VGND VGND VPWR VPWR registers\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31989_ clknet_leaf_22_CLK _00160_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_252_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_252_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24530_ _09598_ registers\[56\]\[40\] _10484_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__mux2_1
X_33728_ clknet_leaf_257_CLK _01842_ VGND VGND VPWR VPWR registers\[41\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_21742_ registers\[0\]\[30\] registers\[1\]\[30\] registers\[2\]\[30\] registers\[3\]\[30\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__mux4_1
XFILLER_240_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24461_ _10448_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
X_33659_ clknet_leaf_277_CLK _01773_ VGND VGND VPWR VPWR registers\[42\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_21673_ registers\[12\]\[28\] registers\[13\]\[28\] registers\[14\]\[28\] registers\[15\]\[28\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__mux4_1
XFILLER_52_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_225_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23412_ _09860_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
X_26200_ _10785_ registers\[44\]\[26\] _11394_ VGND VGND VPWR VPWR _11401_ sky130_fd_sc_hd__mux2_1
X_20624_ _07313_ _07318_ _07321_ _07322_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__a22o_1
X_27180_ _11948_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_1
X_24392_ registers\[57\]\[47\] _10403_ _10389_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__mux2_1
XFILLER_138_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26131_ _11364_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
X_35329_ clknet_leaf_222_CLK _03443_ VGND VGND VPWR VPWR registers\[16\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_23343_ registers\[9\]\[62\] _09823_ _09708_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__mux2_1
XFILLER_71_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20555_ registers\[60\]\[63\] registers\[61\]\[63\] registers\[62\]\[63\] registers\[63\]\[63\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__mux4_1
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26062_ _11328_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
X_23274_ net36 VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__buf_4
X_20486_ registers\[32\]\[61\] registers\[33\]\[61\] registers\[34\]\[61\] registers\[35\]\[61\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__mux4_1
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25013_ net62 VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__buf_4
X_22225_ _07314_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__buf_6
XFILLER_69_1163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_1455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29821_ _13369_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__clkbuf_1
XTAP_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22156_ registers\[44\]\[42\] registers\[45\]\[42\] registers\[46\]\[42\] registers\[47\]\[42\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__mux4_1
XTAP_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1609 _14974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21107_ _07648_ _07792_ _07793_ _07652_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__a22o_1
XFILLER_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29752_ registers\[1\]\[46\] _13031_ _13326_ VGND VGND VPWR VPWR _13333_ sky130_fd_sc_hd__mux2_1
XFILLER_105_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26964_ _11825_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__clkbuf_1
X_22087_ registers\[52\]\[40\] registers\[53\]\[40\] registers\[54\]\[40\] registers\[55\]\[40\]
+ _08605_ _08606_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__mux4_1
XTAP_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28703_ _11788_ registers\[26\]\[28\] _12741_ VGND VGND VPWR VPWR _12750_ sky130_fd_sc_hd__mux2_1
X_25915_ _10770_ registers\[46\]\[19\] _11241_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__mux2_1
X_21038_ registers\[12\]\[10\] registers\[13\]\[10\] registers\[14\]\[10\] registers\[15\]\[10\]
+ _07487_ _07488_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__mux4_1
X_29683_ registers\[1\]\[13\] _12962_ _13293_ VGND VGND VPWR VPWR _13297_ sky130_fd_sc_hd__mux2_1
XFILLER_248_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26895_ _11778_ registers\[3\]\[23\] _11772_ VGND VGND VPWR VPWR _11779_ sky130_fd_sc_hd__mux2_1
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_219_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_491_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_491_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28634_ _12713_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__clkbuf_1
X_25846_ _10835_ registers\[47\]\[50\] _11214_ VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__mux2_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28565_ _12677_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__clkbuf_1
X_25777_ _11178_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
X_22989_ _09588_ registers\[62\]\[35\] _09578_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__mux2_1
XFILLER_43_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_243_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_243_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27516_ _11818_ registers\[35\]\[42\] _12122_ VGND VGND VPWR VPWR _12125_ sky130_fd_sc_hd__mux2_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24728_ _10591_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_1437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28496_ _11851_ registers\[28\]\[58\] _12632_ VGND VGND VPWR VPWR _12641_ sky130_fd_sc_hd__mux2_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27447_ _12088_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__clkbuf_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _09590_ registers\[55\]\[36\] _10547_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__mux2_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17200_ _14500_ VGND VGND VPWR VPWR _15682_ sky130_fd_sc_hd__buf_2
XFILLER_169_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ registers\[20\]\[60\] registers\[21\]\[60\] registers\[22\]\[60\] registers\[23\]\[60\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__mux4_1
XFILLER_204_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27378_ _12052_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17131_ registers\[48\]\[30\] registers\[49\]\[30\] registers\[50\]\[30\] registers\[51\]\[30\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15615_ sky130_fd_sc_hd__mux4_1
X_29117_ net14 VGND VGND VPWR VPWR _12979_ sky130_fd_sc_hd__clkbuf_4
XFILLER_141_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26329_ _10779_ registers\[43\]\[23\] _11465_ VGND VGND VPWR VPWR _11469_ sky130_fd_sc_hd__mux2_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29048_ net1 VGND VGND VPWR VPWR _12931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17062_ _15541_ _15543_ _15546_ _15547_ VGND VGND VPWR VPWR _15548_ sky130_fd_sc_hd__a22o_1
XFILLER_221_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16013_ _14489_ VGND VGND VPWR VPWR _14527_ sky130_fd_sc_hd__buf_12
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31010_ _13995_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _04632_ _04736_ _04737_ _04635_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a22o_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19703_ _06226_ _06426_ _06427_ _06231_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__a22o_1
X_16915_ registers\[44\]\[24\] registers\[45\]\[24\] registers\[46\]\[24\] registers\[47\]\[24\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15405_ sky130_fd_sc_hd__mux4_1
X_32961_ clknet_leaf_294_CLK _01075_ VGND VGND VPWR VPWR registers\[53\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17895_ registers\[28\]\[51\] registers\[29\]\[51\] registers\[30\]\[51\] registers\[31\]\[51\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_482_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_482_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34700_ clknet_leaf_148_CLK _02814_ VGND VGND VPWR VPWR registers\[26\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_31912_ _14469_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19634_ registers\[44\]\[36\] registers\[45\]\[36\] registers\[46\]\[36\] registers\[47\]\[36\]
+ _06156_ _06157_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__mux4_1
X_35680_ clknet_leaf_489_CLK _03794_ VGND VGND VPWR VPWR registers\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16846_ registers\[32\]\[22\] registers\[33\]\[22\] registers\[34\]\[22\] registers\[35\]\[22\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15338_ sky130_fd_sc_hd__mux4_1
X_32892_ clknet_leaf_292_CLK _01006_ VGND VGND VPWR VPWR registers\[54\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_34631_ clknet_leaf_219_CLK _02745_ VGND VGND VPWR VPWR registers\[27\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31843_ _14433_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__clkbuf_1
X_19565_ registers\[40\]\[34\] registers\[41\]\[34\] registers\[42\]\[34\] registers\[43\]\[34\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux4_1
XFILLER_230_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16777_ registers\[56\]\[20\] registers\[57\]\[20\] registers\[58\]\[20\] registers\[59\]\[20\]
+ _15066_ _15199_ VGND VGND VPWR VPWR _15271_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_234_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_234_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18516_ _05077_ _05273_ _05274_ _05086_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__a22o_1
X_34562_ clknet_leaf_229_CLK _02676_ VGND VGND VPWR VPWR registers\[28\]\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31774_ registers\[59\]\[44\] net39 _14392_ VGND VGND VPWR VPWR _14397_ sky130_fd_sc_hd__mux2_1
X_19496_ _05042_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__buf_4
XFILLER_234_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33513_ clknet_leaf_60_CLK _01627_ VGND VGND VPWR VPWR registers\[44\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_18447_ _05204_ _05205_ _05206_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a22o_1
X_30725_ registers\[12\]\[59\] _13058_ _13835_ VGND VGND VPWR VPWR _13845_ sky130_fd_sc_hd__mux2_1
XFILLER_222_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34493_ clknet_leaf_299_CLK _02607_ VGND VGND VPWR VPWR registers\[2\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36232_ clknet_leaf_121_CLK _00117_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dfxtp_1
X_33444_ clknet_leaf_62_CLK _01558_ VGND VGND VPWR VPWR registers\[45\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_18378_ _05078_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__buf_12
X_30656_ registers\[12\]\[26\] _12989_ _13802_ VGND VGND VPWR VPWR _13809_ sky130_fd_sc_hd__mux2_1
XFILLER_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36163_ clknet_leaf_259_CLK _04277_ VGND VGND VPWR VPWR registers\[49\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17329_ _15784_ _15791_ _15800_ _15807_ VGND VGND VPWR VPWR _15808_ sky130_fd_sc_hd__or4_4
X_33375_ clknet_leaf_34_CLK _01489_ VGND VGND VPWR VPWR registers\[46\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_30587_ _13772_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_965 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35114_ clknet_leaf_458_CLK _03228_ VGND VGND VPWR VPWR registers\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32326_ clknet_leaf_154_CLK _00440_ VGND VGND VPWR VPWR registers\[19\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20340_ _06919_ _07045_ _07046_ _06922_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__a22o_1
X_36094_ clknet_leaf_291_CLK _04208_ VGND VGND VPWR VPWR registers\[59\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_49__f_CLK clknet_5_24_0_CLK VGND VGND VPWR VPWR clknet_6_49__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_35045_ clknet_leaf_448_CLK _03159_ VGND VGND VPWR VPWR registers\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_20271_ registers\[40\]\[54\] registers\[41\]\[54\] registers\[42\]\[54\] registers\[43\]\[54\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__mux4_1
X_32257_ clknet_leaf_260_CLK _00371_ VGND VGND VPWR VPWR registers\[39\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22010_ registers\[56\]\[38\] registers\[57\]\[38\] registers\[58\]\[38\] registers\[59\]\[38\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__mux4_1
X_31208_ _14099_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32188_ clknet_leaf_465_CLK _00302_ VGND VGND VPWR VPWR registers\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31139_ _14062_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__clkbuf_1
XTAP_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_233_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23961_ _10153_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35947_ clknet_leaf_400_CLK _04061_ VGND VGND VPWR VPWR registers\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25700_ registers\[48\]\[46\] _10401_ _11130_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_473_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_473_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_22912_ _09535_ registers\[62\]\[10\] _09536_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__mux2_1
XFILLER_57_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26680_ _11653_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__clkbuf_1
X_23892_ _10117_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
X_35878_ clknet_leaf_463_CLK _03992_ VGND VGND VPWR VPWR registers\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_879 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22843_ _09458_ _09465_ _09472_ _09479_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__or4_4
X_25631_ registers\[48\]\[13\] _10332_ _11097_ VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__mux2_1
X_34829_ clknet_leaf_149_CLK _02943_ VGND VGND VPWR VPWR registers\[24\]\[63\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_225_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_225_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28350_ _12564_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__clkbuf_1
X_22774_ _07296_ _09411_ _09412_ _07302_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__a22o_1
X_25562_ registers\[4\]\[46\] _10401_ _11056_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27301_ registers\[36\]\[4\] _10313_ _12007_ VGND VGND VPWR VPWR _12012_ sky130_fd_sc_hd__mux2_1
X_24513_ _09582_ registers\[56\]\[32\] _10473_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__mux2_1
X_21725_ registers\[44\]\[30\] registers\[45\]\[30\] registers\[46\]\[30\] registers\[47\]\[30\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__mux4_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28281_ _12505_ VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__buf_4
XFILLER_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25493_ registers\[4\]\[13\] _10332_ _11023_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__mux2_1
XFILLER_223_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27232_ _11975_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24444_ _10438_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__buf_12
XFILLER_205_1432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21656_ _07316_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__buf_6
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20607_ _07305_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__buf_4
XFILLER_21_971 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27163_ _11939_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__clkbuf_1
X_24375_ _10392_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21587_ _07983_ _08258_ _08259_ _07989_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__a22o_1
XFILLER_193_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26114_ _11355_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
X_23326_ _09812_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
X_20538_ _05107_ _07237_ _07238_ _05117_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__a22o_1
X_27094_ _11801_ registers\[38\]\[34\] _11898_ VGND VGND VPWR VPWR _11903_ sky130_fd_sc_hd__mux2_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23257_ registers\[9\]\[36\] _09766_ _09754_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__mux2_1
X_26045_ _11319_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
X_20469_ registers\[8\]\[60\] registers\[9\]\[60\] registers\[10\]\[60\] registers\[11\]\[60\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__mux4_1
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22208_ _08858_ _08863_ _08759_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__o21ba_1
XTAP_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23188_ _09724_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
XTAP_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1406 _00177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29804_ _13360_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_234_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1417 _00182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22139_ registers\[24\]\[41\] registers\[25\]\[41\] registers\[26\]\[41\] registers\[27\]\[41\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__mux4_1
XFILLER_239_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1428 _04921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27996_ _12378_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1439 _05059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_960 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29735_ registers\[1\]\[38\] _13014_ _13315_ VGND VGND VPWR VPWR _13324_ sky130_fd_sc_hd__mux2_1
XTAP_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26947_ _11729_ VGND VGND VPWR VPWR _11814_ sky130_fd_sc_hd__buf_4
XFILLER_43_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_464_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_464_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16700_ _14998_ _15194_ _15195_ _15001_ VGND VGND VPWR VPWR _15196_ sky130_fd_sc_hd__a22o_1
XFILLER_248_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29666_ registers\[1\]\[5\] _12945_ _13282_ VGND VGND VPWR VPWR _13288_ sky130_fd_sc_hd__mux2_1
X_17680_ _04294_ _04460_ _04461_ _04299_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a22o_1
XTAP_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26878_ net10 VGND VGND VPWR VPWR _11767_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28617_ _11837_ registers\[27\]\[51\] _12703_ VGND VGND VPWR VPWR _12705_ sky130_fd_sc_hd__mux2_1
X_16631_ _15125_ _15128_ _14926_ VGND VGND VPWR VPWR _15129_ sky130_fd_sc_hd__o21ba_1
X_25829_ _10819_ registers\[47\]\[42\] _11203_ VGND VGND VPWR VPWR _11206_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29597_ _13251_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_216_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_216_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19350_ _05883_ _06083_ _06084_ _05888_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__a22o_1
X_16562_ registers\[44\]\[14\] registers\[45\]\[14\] registers\[46\]\[14\] registers\[47\]\[14\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _15062_ sky130_fd_sc_hd__mux4_1
X_28548_ _12668_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18301_ net80 net79 VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__nor2b_4
XFILLER_245_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19281_ registers\[44\]\[26\] registers\[45\]\[26\] registers\[46\]\[26\] registers\[47\]\[26\]
+ _05813_ _05814_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__mux4_1
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28479_ _12576_ VGND VGND VPWR VPWR _12632_ sky130_fd_sc_hd__buf_4
X_16493_ registers\[32\]\[12\] registers\[33\]\[12\] registers\[34\]\[12\] registers\[35\]\[12\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _14995_ sky130_fd_sc_hd__mux4_1
XFILLER_245_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18232_ registers\[12\]\[62\] registers\[13\]\[62\] registers\[14\]\[62\] registers\[15\]\[62\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__mux4_1
X_30510_ _13732_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31490_ _14247_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30441_ _09802_ registers\[14\]\[52\] _13693_ VGND VGND VPWR VPWR _13696_ sky130_fd_sc_hd__mux2_1
X_18163_ registers\[48\]\[60\] registers\[49\]\[60\] registers\[50\]\[60\] registers\[51\]\[60\]
+ _14542_ _14607_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__mux4_1
XFILLER_157_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17114_ registers\[28\]\[29\] registers\[29\]\[29\] registers\[30\]\[29\] registers\[31\]\[29\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15599_ sky130_fd_sc_hd__mux4_1
X_33160_ clknet_leaf_192_CLK _01274_ VGND VGND VPWR VPWR registers\[50\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18094_ _04863_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_2
X_30372_ _13659_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_209_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_946 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32111_ clknet_leaf_468_CLK _00026_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dfxtp_1
XFILLER_143_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17045_ _15528_ _15531_ _15302_ VGND VGND VPWR VPWR _15532_ sky130_fd_sc_hd__o21ba_1
X_33091_ clknet_leaf_270_CLK _01205_ VGND VGND VPWR VPWR registers\[51\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32042_ clknet_leaf_408_CLK _00220_ VGND VGND VPWR VPWR registers\[62\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ registers\[32\]\[18\] registers\[33\]\[18\] registers\[34\]\[18\] registers\[35\]\[18\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__mux4_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35801_ clknet_leaf_14_CLK _03915_ VGND VGND VPWR VPWR registers\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_17947_ registers\[48\]\[53\] registers\[49\]\[53\] registers\[50\]\[53\] registers\[51\]\[53\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__mux4_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33993_ clknet_leaf_261_CLK _02107_ VGND VGND VPWR VPWR registers\[37\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_455_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_455_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_239_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35732_ clknet_leaf_80_CLK _03846_ VGND VGND VPWR VPWR registers\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_32944_ clknet_leaf_368_CLK _01058_ VGND VGND VPWR VPWR registers\[53\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_17878_ registers\[56\]\[51\] registers\[57\]\[51\] registers\[58\]\[51\] registers\[59\]\[51\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux4_1
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19617_ _06031_ _06343_ _06344_ _06034_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__a22o_1
X_16829_ registers\[12\]\[21\] registers\[13\]\[21\] registers\[14\]\[21\] registers\[15\]\[21\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15322_ sky130_fd_sc_hd__mux4_1
XFILLER_54_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35663_ clknet_leaf_135_CLK _03777_ VGND VGND VPWR VPWR registers\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32875_ clknet_leaf_422_CLK _00989_ VGND VGND VPWR VPWR registers\[54\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_207_CLK clknet_6_52__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_207_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_207_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31826_ _14424_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__clkbuf_1
X_19548_ registers\[0\]\[33\] registers\[1\]\[33\] registers\[2\]\[33\] registers\[3\]\[33\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux4_1
X_34614_ clknet_leaf_312_CLK _02728_ VGND VGND VPWR VPWR registers\[27\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_35594_ clknet_leaf_157_CLK _03708_ VGND VGND VPWR VPWR registers\[12\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_222_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34545_ clknet_leaf_385_CLK _02659_ VGND VGND VPWR VPWR registers\[28\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_19479_ registers\[8\]\[31\] registers\[9\]\[31\] registers\[10\]\[31\] registers\[11\]\[31\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__mux4_1
X_31757_ registers\[59\]\[36\] net30 _14381_ VGND VGND VPWR VPWR _14388_ sky130_fd_sc_hd__mux2_1
XFILLER_55_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21510_ _08162_ _08169_ _08178_ _08185_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__or4_4
X_30708_ _13836_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22490_ _08958_ _09136_ _09137_ _08961_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__a22o_1
X_34476_ clknet_leaf_388_CLK _02590_ VGND VGND VPWR VPWR registers\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_31688_ registers\[59\]\[3\] net34 _14348_ VGND VGND VPWR VPWR _14352_ sky130_fd_sc_hd__mux2_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1089 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33427_ clknet_leaf_129_CLK _01541_ VGND VGND VPWR VPWR registers\[45\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_36215_ clknet_leaf_115_CLK _00099_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dfxtp_1
X_21441_ _08118_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30639_ registers\[12\]\[18\] _12972_ _13791_ VGND VGND VPWR VPWR _13800_ sky130_fd_sc_hd__mux2_1
XFILLER_147_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36146_ clknet_leaf_365_CLK _04260_ VGND VGND VPWR VPWR registers\[49\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_24160_ _10259_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
X_33358_ clknet_leaf_130_CLK _01472_ VGND VGND VPWR VPWR registers\[46\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21372_ registers\[44\]\[20\] registers\[45\]\[20\] registers\[46\]\[20\] registers\[47\]\[20\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__mux4_2
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23111_ net63 VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__buf_4
X_20323_ registers\[4\]\[55\] registers\[5\]\[55\] registers\[6\]\[55\] registers\[7\]\[55\]
+ _06795_ _06796_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__mux4_1
X_32309_ clknet_leaf_416_CLK _00423_ VGND VGND VPWR VPWR registers\[19\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_24091_ _10222_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_1
X_36077_ clknet_leaf_372_CLK _04191_ VGND VGND VPWR VPWR registers\[59\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_33289_ clknet_leaf_208_CLK _01403_ VGND VGND VPWR VPWR registers\[48\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23042_ _09624_ registers\[62\]\[52\] _09620_ VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__mux2_1
X_35028_ clknet_leaf_98_CLK _03142_ VGND VGND VPWR VPWR registers\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_20254_ registers\[0\]\[53\] registers\[1\]\[53\] registers\[2\]\[53\] registers\[3\]\[53\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__mux4_1
XFILLER_190_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27850_ _12301_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20185_ registers\[8\]\[51\] registers\[9\]\[51\] registers\[10\]\[51\] registers\[11\]\[51\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__mux4_1
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_854 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26801_ registers\[40\]\[54\] _10418_ _11713_ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__mux2_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27781_ registers\[33\]\[39\] _10386_ _12255_ VGND VGND VPWR VPWR _12265_ sky130_fd_sc_hd__mux2_1
X_24993_ _10728_ registers\[52\]\[0\] _10731_ VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__mux2_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29520_ _13210_ VGND VGND VPWR VPWR _13211_ sky130_fd_sc_hd__buf_4
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_446_CLK clknet_6_9__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_446_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_218_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26732_ registers\[40\]\[21\] _10349_ _11680_ VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__mux2_1
X_23944_ _09619_ registers\[60\]\[50\] _10144_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__mux2_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29451_ _09756_ registers\[21\]\[31\] _13173_ VGND VGND VPWR VPWR _13175_ sky130_fd_sc_hd__mux2_1
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26663_ _10842_ registers\[41\]\[53\] _11641_ VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__mux2_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_804 _08973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _10108_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_815 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_28402_ _11757_ registers\[28\]\[13\] _12588_ VGND VGND VPWR VPWR _12592_ sky130_fd_sc_hd__mux2_1
XANTENNA_826 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25614_ registers\[48\]\[5\] _10315_ _11086_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__mux2_1
XANTENNA_837 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29382_ _09825_ registers\[22\]\[63\] _13068_ VGND VGND VPWR VPWR _13138_ sky130_fd_sc_hd__mux2_1
X_22826_ registers\[52\]\[62\] registers\[53\]\[62\] registers\[54\]\[62\] registers\[55\]\[62\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__mux4_1
XFILLER_44_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_848 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26594_ _10772_ registers\[41\]\[20\] _11608_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__mux2_1
XANTENNA_859 _09277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_819 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28333_ _12555_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25545_ registers\[4\]\[38\] _10384_ _11045_ VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__mux2_1
X_22757_ _09148_ _09394_ _09395_ _09153_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__a22o_1
XFILLER_164_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21708_ registers\[4\]\[29\] registers\[5\]\[29\] registers\[6\]\[29\] registers\[7\]\[29\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__mux4_1
X_28264_ _12519_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__clkbuf_1
X_22688_ _09104_ _09328_ _09329_ _09107_ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__a22o_1
XFILLER_212_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25476_ registers\[4\]\[5\] _10315_ _11012_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__mux2_1
XFILLER_200_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_858 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27215_ _11966_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24427_ _10427_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
X_21639_ registers\[24\]\[27\] registers\[25\]\[27\] registers\[26\]\[27\] registers\[27\]\[27\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__mux4_1
X_28195_ _11820_ registers\[30\]\[43\] _12479_ VGND VGND VPWR VPWR _12483_ sky130_fd_sc_hd__mux2_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27146_ _11853_ registers\[38\]\[59\] _11920_ VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__mux2_1
XFILLER_126_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24358_ registers\[57\]\[36\] _10380_ _10368_ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__mux2_1
XFILLER_126_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23309_ _09801_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24289_ net6 VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__clkbuf_8
X_27077_ _11784_ registers\[38\]\[26\] _11887_ VGND VGND VPWR VPWR _11894_ sky130_fd_sc_hd__mux2_1
XFILLER_181_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26028_ _11310_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_6_32__f_CLK clknet_5_16_0_CLK VGND VGND VPWR VPWR clknet_6_32__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1203 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18850_ registers\[24\]\[13\] registers\[25\]\[13\] registers\[26\]\[13\] registers\[27\]\[13\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__mux4_1
XTAP_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1214 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1225 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17801_ _04340_ _04577_ _04578_ _04343_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__a22o_1
XFILLER_136_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1236 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1247 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1258 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18781_ registers\[16\]\[11\] registers\[17\]\[11\] registers\[18\]\[11\] registers\[19\]\[11\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__mux4_1
X_15993_ _14491_ _14498_ _14501_ _14506_ VGND VGND VPWR VPWR _14507_ sky130_fd_sc_hd__a22o_1
XTAP_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27979_ _12369_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1269 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_437_CLK clknet_6_14__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_437_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_236_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ registers\[48\]\[47\] registers\[49\]\[47\] registers\[50\]\[47\] registers\[51\]\[47\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__mux4_1
X_29718_ _13281_ VGND VGND VPWR VPWR _13315_ sky130_fd_sc_hd__buf_4
XTAP_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30990_ _13984_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__clkbuf_1
XTAP_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29649_ _13278_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__clkbuf_1
X_17663_ registers\[52\]\[45\] registers\[53\]\[45\] registers\[54\]\[45\] registers\[55\]\[45\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__mux4_1
XFILLER_169_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19402_ _06098_ _06134_ _06135_ _06102_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__a22o_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _14801_ _15111_ _15112_ _14804_ VGND VGND VPWR VPWR _15113_ sky130_fd_sc_hd__a22o_1
X_32660_ clknet_leaf_69_CLK _00774_ VGND VGND VPWR VPWR registers\[57\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17594_ registers\[48\]\[43\] registers\[49\]\[43\] registers\[50\]\[43\] registers\[51\]\[43\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__mux4_1
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19333_ registers\[0\]\[27\] registers\[1\]\[27\] registers\[2\]\[27\] registers\[3\]\[27\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__mux4_1
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31611_ _14311_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16545_ _14520_ VGND VGND VPWR VPWR _15046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32591_ clknet_leaf_173_CLK _00705_ VGND VGND VPWR VPWR registers\[58\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34330_ clknet_leaf_4_CLK _02444_ VGND VGND VPWR VPWR registers\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31542_ _14274_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19264_ _05688_ _06000_ _06001_ _05691_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__a22o_1
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16476_ registers\[12\]\[11\] registers\[13\]\[11\] registers\[14\]\[11\] registers\[15\]\[11\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14979_ sky130_fd_sc_hd__mux4_1
XFILLER_148_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18215_ registers\[40\]\[62\] registers\[41\]\[62\] registers\[42\]\[62\] registers\[43\]\[62\]
+ _14534_ _14535_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__mux4_1
X_34261_ clknet_leaf_121_CLK _02375_ VGND VGND VPWR VPWR registers\[32\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_31473_ _14238_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__clkbuf_1
X_19195_ registers\[0\]\[23\] registers\[1\]\[23\] registers\[2\]\[23\] registers\[3\]\[23\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__mux4_1
XFILLER_12_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36000_ clknet_leaf_444_CLK _04114_ VGND VGND VPWR VPWR registers\[63\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_33212_ clknet_leaf_299_CLK _01326_ VGND VGND VPWR VPWR registers\[4\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18146_ registers\[24\]\[59\] registers\[25\]\[59\] registers\[26\]\[59\] registers\[27\]\[59\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__mux4_1
X_30424_ _09784_ registers\[14\]\[44\] _13682_ VGND VGND VPWR VPWR _13687_ sky130_fd_sc_hd__mux2_1
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34192_ clknet_leaf_128_CLK _02306_ VGND VGND VPWR VPWR registers\[33\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33143_ clknet_leaf_335_CLK _01257_ VGND VGND VPWR VPWR registers\[50\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_18077_ _04548_ _04845_ _04846_ _04552_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a22o_1
XFILLER_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30355_ _09681_ registers\[14\]\[11\] _13649_ VGND VGND VPWR VPWR _13651_ sky130_fd_sc_hd__mux2_1
XFILLER_116_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_236_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17028_ registers\[60\]\[27\] registers\[61\]\[27\] registers\[62\]\[27\] registers\[63\]\[27\]
+ _15413_ _15207_ VGND VGND VPWR VPWR _15515_ sky130_fd_sc_hd__mux4_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33074_ clknet_leaf_364_CLK _01188_ VGND VGND VPWR VPWR registers\[51\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30286_ registers\[15\]\[43\] _13025_ _13610_ VGND VGND VPWR VPWR _13614_ sky130_fd_sc_hd__mux2_1
XFILLER_125_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32025_ clknet_leaf_66_CLK _00203_ VGND VGND VPWR VPWR registers\[62\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ registers\[8\]\[17\] registers\[9\]\[17\] registers\[10\]\[17\] registers\[11\]\[17\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__mux4_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1770 _09666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_428_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_428_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1781 _12718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21990_ _08615_ _08650_ _08651_ _08618_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__a22o_1
X_33976_ clknet_leaf_337_CLK _02090_ VGND VGND VPWR VPWR registers\[37\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_1377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35715_ clknet_leaf_241_CLK _03829_ VGND VGND VPWR VPWR registers\[10\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_20941_ _07632_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
X_32927_ clknet_leaf_46_CLK _01041_ VGND VGND VPWR VPWR registers\[53\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20872_ registers\[40\]\[6\] registers\[41\]\[6\] registers\[42\]\[6\] registers\[43\]\[6\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__mux4_1
XFILLER_198_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35646_ clknet_leaf_295_CLK _03760_ VGND VGND VPWR VPWR registers\[11\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_23660_ _09993_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32858_ clknet_leaf_67_CLK _00972_ VGND VGND VPWR VPWR registers\[54\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22611_ _09251_ _09254_ _09083_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__o21ba_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31809_ registers\[59\]\[61\] net58 _14347_ VGND VGND VPWR VPWR _14415_ sky130_fd_sc_hd__mux2_1
X_23591_ _09957_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
X_32789_ clknet_leaf_182_CLK _00903_ VGND VGND VPWR VPWR registers\[55\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_35577_ clknet_leaf_303_CLK _03691_ VGND VGND VPWR VPWR registers\[12\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22542_ registers\[44\]\[53\] registers\[45\]\[53\] registers\[46\]\[53\] registers\[47\]\[53\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__mux4_1
X_25330_ _10939_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__clkbuf_1
X_34528_ clknet_leaf_488_CLK _02642_ VGND VGND VPWR VPWR registers\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22473_ _08805_ _09119_ _09120_ _08810_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__a22o_1
X_25261_ _10902_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34459_ clknet_leaf_478_CLK _02573_ VGND VGND VPWR VPWR registers\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_27000_ _11849_ registers\[3\]\[57\] _11835_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__mux2_1
X_24212_ _10286_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_21424_ _07991_ _08100_ _08101_ _07995_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__a22o_1
X_25192_ _10866_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24143_ _10250_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
X_21355_ registers\[4\]\[19\] registers\[5\]\[19\] registers\[6\]\[19\] registers\[7\]\[19\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__mux4_1
X_36129_ clknet_leaf_42_CLK _04243_ VGND VGND VPWR VPWR registers\[49\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20306_ registers\[32\]\[55\] registers\[33\]\[55\] registers\[34\]\[55\] registers\[35\]\[55\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__mux4_1
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24074_ _10213_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__clkbuf_1
X_28951_ _12880_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21286_ registers\[24\]\[17\] registers\[25\]\[17\] registers\[26\]\[17\] registers\[27\]\[17\]
+ _07867_ _07868_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__mux4_1
XFILLER_162_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23025_ net42 VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__clkbuf_4
X_27902_ registers\[32\]\[32\] _10372_ _12326_ VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__mux2_1
X_20237_ _06924_ _06931_ _06938_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__or4_4
XFILLER_104_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28882_ _11832_ registers\[25\]\[49\] _12834_ VGND VGND VPWR VPWR _12844_ sky130_fd_sc_hd__mux2_1
XFILLER_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27833_ _09653_ _11084_ VGND VGND VPWR VPWR _12292_ sky130_fd_sc_hd__nor2_8
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20168_ _06872_ _06879_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__o21ba_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_419_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_419_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27764_ _12256_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__clkbuf_1
X_24976_ _10721_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__clkbuf_1
X_20099_ registers\[44\]\[49\] registers\[45\]\[49\] registers\[46\]\[49\] registers\[47\]\[49\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__mux4_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29503_ _09810_ registers\[21\]\[56\] _13195_ VGND VGND VPWR VPWR _13202_ sky130_fd_sc_hd__mux2_1
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26715_ registers\[40\]\[13\] _10332_ _11669_ VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__mux2_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _09603_ registers\[60\]\[42\] _10133_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__mux2_1
XFILLER_40_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27695_ _12219_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_933 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_601 _05088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_612 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29434_ _09730_ registers\[21\]\[23\] _13162_ VGND VGND VPWR VPWR _13166_ sky130_fd_sc_hd__mux2_1
XANTENNA_623 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26646_ _10825_ registers\[41\]\[45\] _11630_ VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__mux2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_634 _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23858_ _10099_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_645 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_656 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ registers\[28\]\[61\] registers\[29\]\[61\] registers\[30\]\[61\] registers\[31\]\[61\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__mux4_1
X_29365_ _13129_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_667 _05396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_678 _05882_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26577_ _10756_ registers\[41\]\[12\] _11597_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__mux2_1
XFILLER_246_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23789_ _09601_ registers\[29\]\[41\] _10061_ VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__mux2_1
XANTENNA_689 _06473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16330_ registers\[4\]\[7\] registers\[5\]\[7\] registers\[6\]\[7\] registers\[7\]\[7\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14837_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28316_ _12546_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25528_ _11011_ VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__buf_6
XFILLER_185_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29296_ _13093_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_242_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28247_ _12510_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__clkbuf_1
X_16261_ _14570_ _14768_ _14769_ _14582_ VGND VGND VPWR VPWR _14770_ sky130_fd_sc_hd__a22o_1
X_25459_ _11006_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18000_ registers\[20\]\[54\] registers\[21\]\[54\] registers\[22\]\[54\] registers\[23\]\[54\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux4_1
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16192_ _14573_ VGND VGND VPWR VPWR _14703_ sky130_fd_sc_hd__buf_4
X_28178_ _11803_ registers\[30\]\[35\] _12468_ VGND VGND VPWR VPWR _12474_ sky130_fd_sc_hd__mux2_1
XFILLER_12_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27129_ _11921_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30140_ registers\[16\]\[38\] _13014_ _13528_ VGND VGND VPWR VPWR _13537_ sky130_fd_sc_hd__mux2_1
XFILLER_138_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19951_ _06669_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
X_18902_ _05404_ _05648_ _05649_ _05410_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a22o_1
X_30071_ registers\[16\]\[5\] _12945_ _13495_ VGND VGND VPWR VPWR _13501_ sky130_fd_sc_hd__mux2_1
XFILLER_136_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1000 _11820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_19882_ _06530_ _06601_ _06602_ _06535_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__a22o_1
XFILLER_106_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1011 _11935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1022 _12505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1033 _12966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1044 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18833_ _05579_ _05582_ _05475_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__o21ba_1
XTAP_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1055 _13494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1066 _14063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1077 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18764_ _05204_ _05514_ _05515_ _05207_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__a22o_1
X_33830_ clknet_leaf_456_CLK _01944_ VGND VGND VPWR VPWR registers\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1088 _14504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1099 _14527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15976_ _14489_ VGND VGND VPWR VPWR _14490_ sky130_fd_sc_hd__buf_12
XFILLER_23_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _04289_ _04492_ _04495_ _04292_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__a22o_1
XFILLER_76_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33761_ clknet_leaf_39_CLK _01875_ VGND VGND VPWR VPWR registers\[40\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_30973_ _13975_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__clkbuf_1
X_18695_ registers\[52\]\[9\] registers\[53\]\[9\] registers\[54\]\[9\] registers\[55\]\[9\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__mux4_1
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35500_ clknet_leaf_392_CLK _03614_ VGND VGND VPWR VPWR registers\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32712_ clknet_leaf_209_CLK _00826_ VGND VGND VPWR VPWR registers\[57\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_17646_ registers\[28\]\[44\] registers\[29\]\[44\] registers\[30\]\[44\] registers\[31\]\[44\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__mux4_1
XFILLER_97_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33692_ clknet_leaf_27_CLK _01806_ VGND VGND VPWR VPWR registers\[41\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_999 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32643_ clknet_leaf_266_CLK _00757_ VGND VGND VPWR VPWR registers\[58\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_35431_ clknet_leaf_461_CLK _03545_ VGND VGND VPWR VPWR registers\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17577_ _04289_ _04360_ _04361_ _04292_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__a22o_1
XFILLER_51_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19316_ registers\[40\]\[27\] registers\[41\]\[27\] registers\[42\]\[27\] registers\[43\]\[27\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__mux4_1
X_35362_ clknet_leaf_468_CLK _03476_ VGND VGND VPWR VPWR registers\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_16528_ registers\[32\]\[13\] registers\[33\]\[13\] registers\[34\]\[13\] registers\[35\]\[13\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15029_ sky130_fd_sc_hd__mux4_1
XFILLER_189_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32574_ clknet_leaf_197_CLK _00688_ VGND VGND VPWR VPWR registers\[5\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34313_ clknet_leaf_237_CLK _02427_ VGND VGND VPWR VPWR registers\[32\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_31525_ _09806_ registers\[6\]\[54\] _14261_ VGND VGND VPWR VPWR _14266_ sky130_fd_sc_hd__mux2_1
X_19247_ registers\[32\]\[25\] registers\[33\]\[25\] registers\[34\]\[25\] registers\[35\]\[25\]
+ _05780_ _05781_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__mux4_1
X_16459_ registers\[40\]\[11\] registers\[41\]\[11\] registers\[42\]\[11\] registers\[43\]\[11\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14962_ sky130_fd_sc_hd__mux4_1
X_35293_ clknet_leaf_5_CLK _03407_ VGND VGND VPWR VPWR registers\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_34244_ clknet_leaf_246_CLK _02358_ VGND VGND VPWR VPWR registers\[33\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31456_ _09702_ registers\[6\]\[21\] _14228_ VGND VGND VPWR VPWR _14230_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19178_ _05895_ _05902_ _05909_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__or4_4
XFILLER_117_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18129_ registers\[36\]\[59\] registers\[37\]\[59\] registers\[38\]\[59\] registers\[39\]\[59\]
+ _14572_ _14574_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux4_1
X_30407_ _09766_ registers\[14\]\[36\] _13671_ VGND VGND VPWR VPWR _13678_ sky130_fd_sc_hd__mux2_1
X_34175_ clknet_leaf_269_CLK _02289_ VGND VGND VPWR VPWR registers\[34\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_31387_ _14193_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21140_ _07822_ _07825_ _07719_ _07720_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__o211a_1
X_33126_ clknet_leaf_439_CLK _01240_ VGND VGND VPWR VPWR registers\[50\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_30338_ _09664_ registers\[14\]\[3\] _13638_ VGND VGND VPWR VPWR _13642_ sky130_fd_sc_hd__mux2_1
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21071_ _07648_ _07757_ _07758_ _07652_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__a22o_1
XFILLER_63_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33057_ clknet_leaf_42_CLK _01171_ VGND VGND VPWR VPWR registers\[51\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_30269_ registers\[15\]\[35\] _13008_ _13599_ VGND VGND VPWR VPWR _13605_ sky130_fd_sc_hd__mux2_1
XFILLER_67_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20022_ registers\[40\]\[47\] registers\[41\]\[47\] registers\[42\]\[47\] registers\[43\]\[47\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__mux4_1
X_32008_ clknet_leaf_29_CLK _00181_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24830_ _09624_ registers\[54\]\[52\] _10642_ VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24761_ _10608_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
X_33959_ clknet_leaf_431_CLK _02073_ VGND VGND VPWR VPWR registers\[37\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_21973_ _07356_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__buf_4
XFILLER_227_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26500_ _10814_ registers\[42\]\[40\] _11558_ VGND VGND VPWR VPWR _11559_ sky130_fd_sc_hd__mux2_1
X_23712_ _10022_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20924_ _07325_ _07614_ _07615_ _07336_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__a22o_1
X_27480_ _11782_ registers\[35\]\[25\] _12100_ VGND VGND VPWR VPWR _12106_ sky130_fd_sc_hd__mux2_1
XFILLER_242_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24692_ _10571_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26431_ _11522_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__clkbuf_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _07289_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__buf_4
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35629_ clknet_leaf_391_CLK _03743_ VGND VGND VPWR VPWR registers\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23643_ _09984_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29150_ _13001_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26362_ _10812_ registers\[43\]\[39\] _11476_ VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__mux2_1
X_20786_ _07325_ _07480_ _07481_ _07336_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__a22o_1
X_23574_ _09948_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28101_ _11861_ registers\[31\]\[63\] _12363_ VGND VGND VPWR VPWR _12433_ sky130_fd_sc_hd__mux2_1
XFILLER_168_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25313_ _10929_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__clkbuf_1
X_22525_ registers\[4\]\[52\] registers\[5\]\[52\] registers\[6\]\[52\] registers\[7\]\[52\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__mux4_1
X_29081_ _12954_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__clkbuf_1
X_26293_ _10743_ registers\[43\]\[6\] _11443_ VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__mux2_1
XFILLER_194_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28032_ _12363_ VGND VGND VPWR VPWR _12397_ sky130_fd_sc_hd__buf_4
XFILLER_196_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25244_ _10893_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_1
X_22456_ registers\[24\]\[50\] registers\[25\]\[50\] registers\[26\]\[50\] registers\[27\]\[50\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__mux4_1
XFILLER_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21407_ _08080_ _08081_ _08084_ _08085_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__a22o_1
X_25175_ _10854_ registers\[52\]\[59\] _10836_ VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__mux2_1
X_22387_ _08761_ _09036_ _09037_ _08764_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__a22o_1
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24126_ _10241_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__clkbuf_1
X_21338_ registers\[32\]\[19\] registers\[33\]\[19\] registers\[34\]\[19\] registers\[35\]\[19\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__mux4_1
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29983_ _13454_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28934_ _12871_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24057_ _10204_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__clkbuf_1
X_21269_ registers\[36\]\[17\] registers\[37\]\[17\] registers\[38\]\[17\] registers\[39\]\[17\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__mux4_1
XFILLER_235_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23008_ _09601_ registers\[62\]\[41\] _09599_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__mux2_1
XFILLER_150_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28865_ _12835_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27816_ _12283_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__clkbuf_1
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28796_ _11746_ registers\[25\]\[8\] _12790_ VGND VGND VPWR VPWR _12799_ sky130_fd_sc_hd__mux2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27747_ _12247_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__clkbuf_1
X_24959_ _10712_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _14584_ VGND VGND VPWR VPWR _15974_ sky130_fd_sc_hd__buf_2
XFILLER_233_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _05236_ _05239_ _05074_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__o21ba_1
XFILLER_218_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27678_ registers\[34\]\[54\] _10418_ _12206_ VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__mux2_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_420 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_431 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_442 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29417_ _09689_ registers\[21\]\[15\] _13151_ VGND VGND VPWR VPWR _13157_ sky130_fd_sc_hd__mux2_1
X_17431_ _15901_ _15906_ _15631_ VGND VGND VPWR VPWR _15907_ sky130_fd_sc_hd__o21ba_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26629_ _10808_ registers\[41\]\[37\] _11619_ VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__mux2_1
XANTENNA_453 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_464 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_475 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_486 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29348_ _13120_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__clkbuf_1
X_17362_ _15633_ _15836_ _15839_ _15636_ VGND VGND VPWR VPWR _15840_ sky130_fd_sc_hd__a22o_1
XANTENNA_497 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19101_ _05149_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__clkbuf_4
X_16313_ registers\[44\]\[7\] registers\[45\]\[7\] registers\[46\]\[7\] registers\[47\]\[7\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14820_ sky130_fd_sc_hd__mux4_1
XFILLER_202_964 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29279_ _13084_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__clkbuf_1
X_17293_ registers\[28\]\[34\] registers\[29\]\[34\] registers\[30\]\[34\] registers\[31\]\[34\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15773_ sky130_fd_sc_hd__mux4_1
XFILLER_105_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19032_ _05773_ _05776_ _05508_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__o21ba_1
X_31310_ registers\[7\]\[16\] net8 _14146_ VGND VGND VPWR VPWR _14153_ sky130_fd_sc_hd__mux2_1
X_16244_ registers\[36\]\[5\] registers\[37\]\[5\] registers\[38\]\[5\] registers\[39\]\[5\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _14753_ sky130_fd_sc_hd__mux4_1
XFILLER_186_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32290_ clknet_leaf_474_CLK _00404_ VGND VGND VPWR VPWR registers\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1051 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31241_ _14116_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__clkbuf_1
X_16175_ registers\[32\]\[3\] registers\[33\]\[3\] registers\[34\]\[3\] registers\[35\]\[3\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14686_ sky130_fd_sc_hd__mux4_1
XFILLER_177_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR D1[25] sky130_fd_sc_hd__buf_2
Xoutput118 net118 VGND VGND VPWR VPWR D1[35] sky130_fd_sc_hd__buf_2
XFILLER_182_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31172_ _14080_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__clkbuf_1
Xoutput129 net129 VGND VGND VPWR VPWR D1[45] sky130_fd_sc_hd__buf_2
XFILLER_177_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30123_ _13494_ VGND VGND VPWR VPWR _13528_ sky130_fd_sc_hd__buf_4
XFILLER_138_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19934_ registers\[8\]\[44\] registers\[9\]\[44\] registers\[10\]\[44\] registers\[11\]\[44\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__mux4_1
X_35980_ clknet_leaf_144_CLK _04094_ VGND VGND VPWR VPWR registers\[6\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30054_ _13491_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34931_ clknet_leaf_384_CLK _03045_ VGND VGND VPWR VPWR registers\[22\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_19865_ registers\[52\]\[42\] registers\[53\]\[42\] registers\[54\]\[42\] registers\[55\]\[42\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__mux4_1
X_18816_ registers\[24\]\[12\] registers\[25\]\[12\] registers\[26\]\[12\] registers\[27\]\[12\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__mux4_1
XTAP_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34862_ clknet_leaf_394_CLK _02976_ VGND VGND VPWR VPWR registers\[23\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19796_ _06374_ _06515_ _06518_ _06377_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__a22o_1
XFILLER_110_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33813_ clknet_leaf_80_CLK _01927_ VGND VGND VPWR VPWR registers\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18747_ _05496_ _05497_ _05498_ _05499_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__a22o_1
XFILLER_237_872 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34793_ clknet_leaf_452_CLK _02907_ VGND VGND VPWR VPWR registers\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33744_ clknet_leaf_129_CLK _01858_ VGND VGND VPWR VPWR registers\[40\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18678_ _05150_ _05431_ _05432_ _05160_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__a22o_1
XFILLER_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30956_ registers\[10\]\[40\] _13018_ _13966_ VGND VGND VPWR VPWR _13967_ sky130_fd_sc_hd__mux2_1
XFILLER_110_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17629_ _14541_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__buf_6
XFILLER_52_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33675_ clknet_leaf_159_CLK _01789_ VGND VGND VPWR VPWR registers\[42\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_30887_ _13930_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35414_ clknet_leaf_81_CLK _03528_ VGND VGND VPWR VPWR registers\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_20640_ _07338_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__buf_2
X_32626_ clknet_leaf_363_CLK _00740_ VGND VGND VPWR VPWR registers\[58\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20571_ _05119_ _07269_ _07270_ _05131_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__a22o_1
X_35345_ clknet_leaf_107_CLK _03459_ VGND VGND VPWR VPWR registers\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_32557_ clknet_leaf_390_CLK _00671_ VGND VGND VPWR VPWR registers\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1074 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22310_ _08957_ _08962_ _08759_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__o21ba_1
X_31508_ _09788_ registers\[6\]\[46\] _14250_ VGND VGND VPWR VPWR _14257_ sky130_fd_sc_hd__mux2_1
X_23290_ registers\[9\]\[46\] _09788_ _09776_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__mux2_1
X_35276_ clknet_leaf_147_CLK _03390_ VGND VGND VPWR VPWR registers\[17\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32488_ clknet_leaf_436_CLK _00602_ VGND VGND VPWR VPWR registers\[60\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22241_ _07347_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__buf_6
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31439_ _09685_ registers\[6\]\[13\] _14217_ VGND VGND VPWR VPWR _14221_ sky130_fd_sc_hd__mux2_1
X_34227_ clknet_leaf_349_CLK _02341_ VGND VGND VPWR VPWR registers\[33\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22172_ registers\[4\]\[42\] registers\[5\]\[42\] registers\[6\]\[42\] registers\[7\]\[42\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__mux4_1
X_34158_ clknet_leaf_352_CLK _02272_ VGND VGND VPWR VPWR registers\[34\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21123_ _07737_ _07808_ _07809_ _07742_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__a22o_1
X_33109_ clknet_leaf_69_CLK _01223_ VGND VGND VPWR VPWR registers\[50\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26980_ _11836_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34089_ clknet_leaf_435_CLK _02203_ VGND VGND VPWR VPWR registers\[35\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25931_ _11259_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
X_21054_ _07737_ _07738_ _07741_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__a22o_1
XFILLER_236_1394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20005_ _05059_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__buf_4
X_28650_ _12722_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__clkbuf_1
X_25862_ _10852_ registers\[47\]\[58\] _11214_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__mux2_1
XFILLER_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27601_ _12170_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1018 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24813_ _09607_ registers\[54\]\[44\] _10631_ VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__mux2_1
X_28581_ _11801_ registers\[27\]\[34\] _12681_ VGND VGND VPWR VPWR _12686_ sky130_fd_sc_hd__mux2_1
X_25793_ _10783_ registers\[47\]\[25\] _11181_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__mux2_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27532_ _12077_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__buf_4
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24744_ _09538_ registers\[54\]\[11\] _10598_ VGND VGND VPWR VPWR _10600_ sky130_fd_sc_hd__mux2_1
XFILLER_227_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21956_ _08615_ _08616_ _08617_ _08618_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__a22o_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20907_ _07596_ _07599_ _07399_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__o21ba_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27463_ _11765_ registers\[35\]\[17\] _12089_ VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__mux2_1
X_24675_ _10562_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21887_ _08548_ _08551_ _08416_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__o21ba_1
XFILLER_215_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29202_ _13036_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26414_ _10935_ _11157_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__nand2_8
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23626_ _09975_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_230_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20838_ _07507_ _07516_ _07523_ _07532_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__or4_2
X_27394_ _12060_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29133_ registers\[23\]\[26\] _12989_ _12977_ VGND VGND VPWR VPWR _12990_ sky130_fd_sc_hd__mux2_1
XFILLER_126_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26345_ _11477_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__clkbuf_1
X_23557_ _09644_ registers\[19\]\[62\] _09869_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__mux2_1
X_20769_ registers\[20\]\[2\] registers\[21\]\[2\] registers\[22\]\[2\] registers\[23\]\[2\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__mux4_1
XFILLER_168_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22508_ _07324_ VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__buf_4
X_29064_ net45 VGND VGND VPWR VPWR _12943_ sky130_fd_sc_hd__buf_2
XFILLER_168_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26276_ _11440_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23488_ _09575_ registers\[19\]\[29\] _09892_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28015_ _12388_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25227_ _10884_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22439_ registers\[60\]\[50\] registers\[61\]\[50\] registers\[62\]\[50\] registers\[63\]\[50\]
+ _08884_ _09021_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__mux4_1
XFILLER_104_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25158_ _10843_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24109_ _10231_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__buf_12
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17980_ registers\[48\]\[54\] registers\[49\]\[54\] registers\[50\]\[54\] registers\[51\]\[54\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__mux4_1
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25089_ _10796_ registers\[52\]\[31\] _10794_ VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__mux2_1
X_29966_ _13445_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16931_ registers\[12\]\[24\] registers\[13\]\[24\] registers\[14\]\[24\] registers\[15\]\[24\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15421_ sky130_fd_sc_hd__mux4_1
XFILLER_46_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28917_ registers\[24\]\[1\] _10307_ _12861_ VGND VGND VPWR VPWR _12863_ sky130_fd_sc_hd__mux2_1
XFILLER_104_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29897_ _13409_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16862_ registers\[8\]\[22\] registers\[9\]\[22\] registers\[10\]\[22\] registers\[11\]\[22\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15354_ sky130_fd_sc_hd__mux4_1
X_19650_ _05116_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__buf_4
X_28848_ _12826_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18601_ _05143_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__buf_4
XFILLER_133_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19581_ registers\[8\]\[34\] registers\[9\]\[34\] registers\[10\]\[34\] registers\[11\]\[34\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__mux4_1
XFILLER_92_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28779_ _12789_ VGND VGND VPWR VPWR _12790_ sky130_fd_sc_hd__clkbuf_8
X_16793_ _15144_ _15285_ _15286_ _15147_ VGND VGND VPWR VPWR _15287_ sky130_fd_sc_hd__a22o_1
XFILLER_237_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18532_ registers\[16\]\[4\] registers\[17\]\[4\] registers\[18\]\[4\] registers\[19\]\[4\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__mux4_1
X_30810_ _09764_ registers\[11\]\[35\] _13884_ VGND VGND VPWR VPWR _13890_ sky130_fd_sc_hd__mux2_1
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31790_ _14405_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__clkbuf_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30741_ _09662_ registers\[11\]\[2\] _13851_ VGND VGND VPWR VPWR _13854_ sky130_fd_sc_hd__mux2_1
X_18463_ registers\[24\]\[2\] registers\[25\]\[2\] registers\[26\]\[2\] registers\[27\]\[2\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__mux4_1
Xclkbuf_5_4_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_4_0_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_248_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_261 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _14500_ VGND VGND VPWR VPWR _15890_ sky130_fd_sc_hd__clkbuf_4
X_33460_ clknet_leaf_345_CLK _01574_ VGND VGND VPWR VPWR registers\[45\]\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _05156_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__buf_4
X_30672_ _13817_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_283 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_294 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32411_ clknet_leaf_1_CLK _00525_ VGND VGND VPWR VPWR registers\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_17345_ _15549_ _15819_ _15822_ _15553_ VGND VGND VPWR VPWR _15823_ sky130_fd_sc_hd__a22o_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33391_ clknet_leaf_362_CLK _01505_ VGND VGND VPWR VPWR registers\[46\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32342_ clknet_leaf_66_CLK _00456_ VGND VGND VPWR VPWR registers\[61\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_35130_ clknet_leaf_302_CLK _03244_ VGND VGND VPWR VPWR registers\[1\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17276_ _14541_ VGND VGND VPWR VPWR _15756_ sky130_fd_sc_hd__buf_6
XFILLER_140_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19015_ _05755_ _05757_ _05758_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__a22o_1
X_16227_ _14570_ _14735_ _14736_ _14582_ VGND VGND VPWR VPWR _14737_ sky130_fd_sc_hd__a22o_1
X_35061_ clknet_leaf_384_CLK _03175_ VGND VGND VPWR VPWR registers\[20\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_32273_ clknet_leaf_101_CLK _00387_ VGND VGND VPWR VPWR registers\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34012_ clknet_leaf_23_CLK _02126_ VGND VGND VPWR VPWR registers\[36\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31224_ _14107_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__clkbuf_1
X_16158_ _14558_ _14668_ _14669_ _14568_ VGND VGND VPWR VPWR _14670_ sky130_fd_sc_hd__a22o_1
XFILLER_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31155_ _14071_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16089_ _14531_ VGND VGND VPWR VPWR _14603_ sky130_fd_sc_hd__buf_12
XFILLER_115_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30106_ _13519_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19917_ _06636_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_35963_ clknet_leaf_304_CLK _04077_ VGND VGND VPWR VPWR registers\[6\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31086_ registers\[0\]\[38\] _13014_ _14026_ VGND VGND VPWR VPWR _14035_ sky130_fd_sc_hd__mux2_1
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30037_ registers\[17\]\[53\] _13046_ _13479_ VGND VGND VPWR VPWR _13483_ sky130_fd_sc_hd__mux2_1
XFILLER_29_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34914_ clknet_leaf_473_CLK _03028_ VGND VGND VPWR VPWR registers\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_19848_ _05076_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35894_ clknet_leaf_319_CLK _04008_ VGND VGND VPWR VPWR registers\[7\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34845_ clknet_leaf_491_CLK _02959_ VGND VGND VPWR VPWR registers\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ registers\[36\]\[40\] registers\[37\]\[40\] registers\[38\]\[40\] registers\[39\]\[40\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__mux4_1
XFILLER_37_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21810_ _08326_ _08475_ _08476_ _08332_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__a22o_1
XFILLER_3_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22790_ _09155_ _09426_ _09427_ _09158_ VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__a22o_1
XFILLER_71_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34776_ clknet_leaf_19_CLK _02890_ VGND VGND VPWR VPWR registers\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31988_ clknet_leaf_22_CLK _00159_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33727_ clknet_leaf_272_CLK _01841_ VGND VGND VPWR VPWR registers\[41\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_21741_ _07349_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__clkbuf_4
X_30939_ registers\[10\]\[32\] _13002_ _13955_ VGND VGND VPWR VPWR _13958_ sky130_fd_sc_hd__mux2_1
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24460_ _09529_ registers\[56\]\[7\] _10440_ VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33658_ clknet_leaf_280_CLK _01772_ VGND VGND VPWR VPWR registers\[42\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_21672_ _08267_ _08341_ _08342_ _08270_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__a22o_1
X_23411_ registers\[39\]\[58\] _09815_ _09851_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__mux2_1
XFILLER_149_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20623_ _07285_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__clkbuf_4
X_32609_ clknet_leaf_43_CLK _00723_ VGND VGND VPWR VPWR registers\[58\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_24391_ net42 VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33589_ clknet_leaf_344_CLK _01703_ VGND VGND VPWR VPWR registers\[43\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_26130_ _10850_ registers\[45\]\[57\] _11356_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35328_ clknet_leaf_222_CLK _03442_ VGND VGND VPWR VPWR registers\[16\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23342_ net59 VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__buf_2
X_20554_ _05136_ _07252_ _07253_ _05146_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__a22o_1
XFILLER_177_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26061_ _10781_ registers\[45\]\[24\] _11323_ VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__mux2_1
X_20485_ registers\[40\]\[61\] registers\[41\]\[61\] registers\[42\]\[61\] registers\[43\]\[61\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__mux4_1
XFILLER_180_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35259_ clknet_leaf_185_CLK _03373_ VGND VGND VPWR VPWR registers\[17\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_23273_ _09777_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25012_ _10744_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22224_ _08875_ _08878_ _08740_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__o21ba_1
XFILLER_146_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22155_ _07324_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__clkbuf_4
X_29820_ registers\[18\]\[14\] _12964_ _13364_ VGND VGND VPWR VPWR _13369_ sky130_fd_sc_hd__mux2_1
XTAP_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21106_ registers\[52\]\[12\] registers\[53\]\[12\] registers\[54\]\[12\] registers\[55\]\[12\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__mux4_1
XFILLER_248_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26963_ _11824_ registers\[3\]\[45\] _11814_ VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__mux2_1
X_29751_ _13332_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__clkbuf_1
X_22086_ registers\[60\]\[40\] registers\[61\]\[40\] registers\[62\]\[40\] registers\[63\]\[40\]
+ _08541_ _08678_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__mux4_1
XTAP_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28702_ _12749_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__clkbuf_1
X_21037_ _07581_ _07722_ _07725_ _07584_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__a22o_1
X_25914_ _11250_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29682_ _13296_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26894_ net16 VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28633_ _11853_ registers\[27\]\[59\] _12703_ VGND VGND VPWR VPWR _12713_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25845_ _11158_ VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__buf_4
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28564_ _11784_ registers\[27\]\[26\] _12670_ VGND VGND VPWR VPWR _12677_ sky130_fd_sc_hd__mux2_1
X_25776_ _10766_ registers\[47\]\[17\] _11170_ VGND VGND VPWR VPWR _11178_ sky130_fd_sc_hd__mux2_1
X_22988_ net29 VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__clkbuf_4
XFILLER_76_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27515_ _12124_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__clkbuf_1
X_24727_ _09521_ registers\[54\]\[3\] _10587_ VGND VGND VPWR VPWR _10591_ sky130_fd_sc_hd__mux2_1
XFILLER_128_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28495_ _12640_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__clkbuf_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21939_ registers\[48\]\[36\] registers\[49\]\[36\] registers\[50\]\[36\] registers\[51\]\[36\]
+ _08329_ _08330_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__mux4_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27446_ _11748_ registers\[35\]\[9\] _12078_ VGND VGND VPWR VPWR _12088_ sky130_fd_sc_hd__mux2_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24658_ _10553_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ registers\[61\]\[21\] _09702_ _09965_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__mux2_1
XFILLER_204_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27377_ registers\[36\]\[40\] _10388_ _12051_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__mux2_1
XFILLER_169_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24589_ _10517_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17130_ registers\[56\]\[30\] registers\[57\]\[30\] registers\[58\]\[30\] registers\[59\]\[30\]
+ _15409_ _15542_ VGND VGND VPWR VPWR _15614_ sky130_fd_sc_hd__mux4_1
X_29116_ _12978_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26328_ _11468_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29047_ _12930_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17061_ _14500_ VGND VGND VPWR VPWR _15547_ sky130_fd_sc_hd__buf_4
X_26259_ _10844_ registers\[44\]\[54\] _11427_ VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__mux2_1
XFILLER_183_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16012_ _14507_ _14523_ _14525_ VGND VGND VPWR VPWR _14526_ sky130_fd_sc_hd__o21ba_1
XFILLER_104_1291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17963_ registers\[16\]\[53\] registers\[17\]\[53\] registers\[18\]\[53\] registers\[19\]\[53\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29949_ registers\[17\]\[11\] _12958_ _13435_ VGND VGND VPWR VPWR _13437_ sky130_fd_sc_hd__mux2_1
X_19702_ registers\[32\]\[38\] registers\[33\]\[38\] registers\[34\]\[38\] registers\[35\]\[38\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16914_ _15334_ _15402_ _15403_ _15339_ VGND VGND VPWR VPWR _15404_ sky130_fd_sc_hd__a22o_1
X_32960_ clknet_leaf_293_CLK _01074_ VGND VGND VPWR VPWR registers\[53\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_17894_ _04632_ _04668_ _04669_ _04635_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__a22o_1
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31911_ _09786_ registers\[49\]\[45\] _14463_ VGND VGND VPWR VPWR _14469_ sky130_fd_sc_hd__mux2_1
X_19633_ _06226_ _06358_ _06359_ _06231_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__a22o_1
XFILLER_238_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16845_ registers\[40\]\[22\] registers\[41\]\[22\] registers\[42\]\[22\] registers\[43\]\[22\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15337_ sky130_fd_sc_hd__mux4_1
X_32891_ clknet_leaf_287_CLK _01005_ VGND VGND VPWR VPWR registers\[54\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34630_ clknet_leaf_218_CLK _02744_ VGND VGND VPWR VPWR registers\[27\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_31842_ _09683_ registers\[49\]\[12\] _14430_ VGND VGND VPWR VPWR _14433_ sky130_fd_sc_hd__mux2_1
X_19564_ _06293_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__buf_2
X_16776_ _15263_ _15268_ _15269_ VGND VGND VPWR VPWR _15270_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18515_ registers\[48\]\[4\] registers\[49\]\[4\] registers\[50\]\[4\] registers\[51\]\[4\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__mux4_1
XFILLER_34_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34561_ clknet_leaf_202_CLK _02675_ VGND VGND VPWR VPWR registers\[28\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_31773_ _14396_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19495_ _05076_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__buf_2
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33512_ clknet_leaf_60_CLK _01626_ VGND VGND VPWR VPWR registers\[44\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_30724_ _13844_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__clkbuf_1
X_18446_ _05130_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__buf_6
X_34492_ clknet_leaf_299_CLK _02606_ VGND VGND VPWR VPWR registers\[2\]\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36231_ clknet_leaf_121_CLK _00116_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dfxtp_1
X_18377_ registers\[24\]\[0\] registers\[25\]\[0\] registers\[26\]\[0\] registers\[27\]\[0\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__mux4_1
XFILLER_159_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33443_ clknet_leaf_58_CLK _01557_ VGND VGND VPWR VPWR registers\[45\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_30655_ _13808_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17328_ _15803_ _15806_ _15645_ VGND VGND VPWR VPWR _15807_ sky130_fd_sc_hd__o21ba_1
XFILLER_239_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36162_ clknet_leaf_263_CLK _04276_ VGND VGND VPWR VPWR registers\[49\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33374_ clknet_leaf_28_CLK _01488_ VGND VGND VPWR VPWR registers\[46\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_30586_ _09813_ registers\[13\]\[57\] _13764_ VGND VGND VPWR VPWR _13772_ sky130_fd_sc_hd__mux2_1
XFILLER_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35113_ clknet_leaf_458_CLK _03227_ VGND VGND VPWR VPWR registers\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_32325_ clknet_leaf_220_CLK _00439_ VGND VGND VPWR VPWR registers\[19\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17259_ registers\[28\]\[33\] registers\[29\]\[33\] registers\[30\]\[33\] registers\[31\]\[33\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15740_ sky130_fd_sc_hd__mux4_1
X_36093_ clknet_leaf_289_CLK _04207_ VGND VGND VPWR VPWR registers\[59\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20270_ _06979_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__buf_4
X_32256_ clknet_leaf_260_CLK _00370_ VGND VGND VPWR VPWR registers\[39\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_35044_ clknet_leaf_472_CLK _03158_ VGND VGND VPWR VPWR registers\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31207_ registers\[8\]\[31\] net25 _14097_ VGND VGND VPWR VPWR _14099_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_170_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_170_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32187_ clknet_leaf_465_CLK _00301_ VGND VGND VPWR VPWR registers\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31138_ registers\[0\]\[63\] _13066_ _13992_ VGND VGND VPWR VPWR _14062_ sky130_fd_sc_hd__mux2_1
XFILLER_130_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23960_ _09636_ registers\[60\]\[58\] _10144_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__mux2_1
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35946_ clknet_leaf_402_CLK _04060_ VGND VGND VPWR VPWR registers\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_31069_ _13992_ VGND VGND VPWR VPWR _14026_ sky130_fd_sc_hd__buf_4
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22911_ _09514_ VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__buf_4
XFILLER_217_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35877_ clknet_leaf_464_CLK _03991_ VGND VGND VPWR VPWR registers\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_23891_ _09567_ registers\[60\]\[25\] _10111_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__mux2_1
X_25630_ _11100_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
X_34828_ clknet_leaf_148_CLK _02942_ VGND VGND VPWR VPWR registers\[24\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_22842_ _09475_ _09478_ _07398_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__o21ba_1
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25561_ _11062_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__clkbuf_1
X_34759_ clknet_leaf_219_CLK _02873_ VGND VGND VPWR VPWR registers\[25\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_22773_ registers\[4\]\[60\] registers\[5\]\[60\] registers\[6\]\[60\] registers\[7\]\[60\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__mux4_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27300_ _12011_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24512_ _10475_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28280_ _12527_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21724_ _07333_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__clkbuf_4
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25492_ _11026_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27231_ _11803_ registers\[37\]\[35\] _11969_ VGND VGND VPWR VPWR _11975_ sky130_fd_sc_hd__mux2_1
XFILLER_240_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24443_ net85 net84 net83 _09512_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__or4b_1
XFILLER_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21655_ _07312_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__buf_4
XFILLER_244_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_240_1335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27162_ _11734_ registers\[37\]\[2\] _11936_ VGND VGND VPWR VPWR _11939_ sky130_fd_sc_hd__mux2_1
X_20606_ _07280_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__buf_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24374_ registers\[57\]\[41\] _10391_ _10389_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__mux2_1
XFILLER_201_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21586_ registers\[48\]\[26\] registers\[49\]\[26\] registers\[50\]\[26\] registers\[51\]\[26\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__mux4_1
X_26113_ _10833_ registers\[45\]\[49\] _11345_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__mux2_1
XFILLER_193_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23325_ registers\[39\]\[27\] _09747_ _09700_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__mux2_1
X_20537_ registers\[16\]\[62\] registers\[17\]\[62\] registers\[18\]\[62\] registers\[19\]\[62\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__mux4_1
X_27093_ _11902_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26044_ _10764_ registers\[45\]\[16\] _11312_ VGND VGND VPWR VPWR _11319_ sky130_fd_sc_hd__mux2_1
X_20468_ _07167_ _07170_ _05102_ _05104_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__o211a_1
X_23256_ net30 VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__buf_2
XFILLER_101_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22207_ _08615_ _08861_ _08862_ _08618_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__a22o_1
XFILLER_10_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_161_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_161_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20399_ registers\[36\]\[58\] registers\[37\]\[58\] registers\[38\]\[58\] registers\[39\]\[58\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__mux4_1
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23187_ registers\[9\]\[11\] _09681_ _09722_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__mux2_1
XTAP_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29803_ registers\[18\]\[6\] _12947_ _13353_ VGND VGND VPWR VPWR _13360_ sky130_fd_sc_hd__mux2_1
XANTENNA_1407 _00177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_234_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1418 _00182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22138_ _08792_ _08795_ _08759_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1429 _04921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27995_ _11755_ registers\[31\]\[12\] _12375_ VGND VGND VPWR VPWR _12378_ sky130_fd_sc_hd__mux2_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29734_ _13323_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26946_ net35 VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__clkbuf_4
XTAP_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22069_ _08423_ _08727_ _08728_ _08428_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__a22o_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29665_ _13287_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__clkbuf_1
X_26877_ _11766_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16630_ _14998_ _15126_ _15127_ _15001_ VGND VGND VPWR VPWR _15128_ sky130_fd_sc_hd__a22o_1
X_28616_ _12704_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__clkbuf_1
X_25828_ _11205_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29596_ registers\[20\]\[36\] _13010_ _13244_ VGND VGND VPWR VPWR _13251_ sky130_fd_sc_hd__mux2_1
XFILLER_62_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16561_ _14991_ _15059_ _15060_ _14996_ VGND VGND VPWR VPWR _15061_ sky130_fd_sc_hd__a22o_1
XFILLER_244_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25759_ _10749_ registers\[47\]\[9\] _11159_ VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__mux2_1
XFILLER_222_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28547_ _11767_ registers\[27\]\[18\] _12659_ VGND VGND VPWR VPWR _12668_ sky130_fd_sc_hd__mux2_1
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18300_ registers\[44\]\[0\] registers\[45\]\[0\] registers\[46\]\[0\] registers\[47\]\[0\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__mux4_1
X_19280_ _05883_ _06015_ _06016_ _05888_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a22o_1
XFILLER_245_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_6_55__f_CLK clknet_5_27_0_CLK VGND VGND VPWR VPWR clknet_6_55__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_28478_ _12631_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__clkbuf_1
X_16492_ registers\[40\]\[12\] registers\[41\]\[12\] registers\[42\]\[12\] registers\[43\]\[12\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _14994_ sky130_fd_sc_hd__mux4_1
XFILLER_231_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18231_ _14491_ _04994_ _04995_ _14501_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__a22o_1
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27429_ _12079_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30440_ _13695_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__clkbuf_1
X_18162_ registers\[56\]\[60\] registers\[57\]\[60\] registers\[58\]\[60\] registers\[59\]\[60\]
+ _04751_ _14603_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__mux4_1
XFILLER_141_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17113_ _15290_ _15596_ _15597_ _15293_ VGND VGND VPWR VPWR _15598_ sky130_fd_sc_hd__a22o_1
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18093_ _04841_ _04848_ _04855_ _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__or4_4
X_30371_ _09697_ registers\[14\]\[19\] _13649_ VGND VGND VPWR VPWR _13659_ sky130_fd_sc_hd__mux2_1
XFILLER_183_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32110_ clknet_leaf_468_CLK _00025_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dfxtp_1
XFILLER_183_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17044_ _15295_ _15529_ _15530_ _15300_ VGND VGND VPWR VPWR _15531_ sky130_fd_sc_hd__a22o_1
X_33090_ clknet_leaf_263_CLK _01204_ VGND VGND VPWR VPWR registers\[51\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32041_ clknet_leaf_451_CLK _00219_ VGND VGND VPWR VPWR registers\[62\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_152_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_152_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ registers\[40\]\[18\] registers\[41\]\[18\] registers\[42\]\[18\] registers\[43\]\[18\]
+ _05541_ _05542_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__mux4_1
XFILLER_174_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35800_ clknet_leaf_14_CLK _03914_ VGND VGND VPWR VPWR registers\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ registers\[56\]\[53\] registers\[57\]\[53\] registers\[58\]\[53\] registers\[59\]\[53\]
+ _04408_ _04541_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__mux4_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33992_ clknet_leaf_237_CLK _02106_ VGND VGND VPWR VPWR registers\[37\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35731_ clknet_leaf_79_CLK _03845_ VGND VGND VPWR VPWR registers\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_32943_ clknet_leaf_368_CLK _01057_ VGND VGND VPWR VPWR registers\[53\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_226_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17877_ _04649_ _04652_ _04611_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__o21ba_1
XFILLER_54_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19616_ registers\[0\]\[35\] registers\[1\]\[35\] registers\[2\]\[35\] registers\[3\]\[35\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__mux4_1
XFILLER_54_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35662_ clknet_leaf_109_CLK _03776_ VGND VGND VPWR VPWR registers\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16828_ _15139_ _15319_ _15320_ _15142_ VGND VGND VPWR VPWR _15321_ sky130_fd_sc_hd__a22o_1
XFILLER_26_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32874_ clknet_leaf_422_CLK _00988_ VGND VGND VPWR VPWR registers\[54\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34613_ clknet_leaf_409_CLK _02727_ VGND VGND VPWR VPWR registers\[27\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_31825_ _09666_ registers\[49\]\[4\] _14419_ VGND VGND VPWR VPWR _14424_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19547_ registers\[8\]\[33\] registers\[9\]\[33\] registers\[10\]\[33\] registers\[11\]\[33\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__mux4_1
X_35593_ clknet_leaf_156_CLK _03707_ VGND VGND VPWR VPWR registers\[12\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_16759_ registers\[16\]\[19\] registers\[17\]\[19\] registers\[18\]\[19\] registers\[19\]\[19\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15254_ sky130_fd_sc_hd__mux4_1
XFILLER_81_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34544_ clknet_leaf_388_CLK _02658_ VGND VGND VPWR VPWR registers\[28\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31756_ _14387_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__clkbuf_1
X_19478_ _06206_ _06209_ _06169_ _06170_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__o211a_1
XFILLER_62_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30707_ registers\[12\]\[50\] _13039_ _13835_ VGND VGND VPWR VPWR _13836_ sky130_fd_sc_hd__mux2_1
X_18429_ _05137_ _05189_ _05190_ _05147_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34475_ clknet_leaf_459_CLK _02589_ VGND VGND VPWR VPWR registers\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31687_ _14351_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36214_ clknet_leaf_115_CLK _00098_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dfxtp_1
X_33426_ clknet_leaf_122_CLK _01540_ VGND VGND VPWR VPWR registers\[45\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21440_ _08096_ _08103_ _08110_ _08117_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__or4_4
X_30638_ _13799_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21371_ _07333_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__clkbuf_4
X_36145_ clknet_leaf_365_CLK _04259_ VGND VGND VPWR VPWR registers\[49\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_33357_ clknet_leaf_172_CLK _01471_ VGND VGND VPWR VPWR registers\[47\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_30569_ _09795_ registers\[13\]\[49\] _13753_ VGND VGND VPWR VPWR _13763_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_391_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_391_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20322_ registers\[12\]\[55\] registers\[13\]\[55\] registers\[14\]\[55\] registers\[15\]\[55\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux4_1
X_23110_ _09673_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_1
X_32308_ clknet_leaf_416_CLK _00422_ VGND VGND VPWR VPWR registers\[19\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_24090_ _09630_ registers\[5\]\[55\] _10216_ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36076_ clknet_leaf_372_CLK _04190_ VGND VGND VPWR VPWR registers\[59\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_33288_ clknet_leaf_208_CLK _01402_ VGND VGND VPWR VPWR registers\[48\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20253_ registers\[8\]\[53\] registers\[9\]\[53\] registers\[10\]\[53\] registers\[11\]\[53\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__mux4_1
X_23041_ net48 VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__buf_4
X_35027_ clknet_leaf_103_CLK _03141_ VGND VGND VPWR VPWR registers\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_143_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_143_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32239_ clknet_leaf_357_CLK _00353_ VGND VGND VPWR VPWR registers\[39\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20184_ _06892_ _06895_ _06855_ _06856_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__o211a_1
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26800_ _11717_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__clkbuf_1
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27780_ _12264_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__clkbuf_1
X_24992_ _10730_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__buf_4
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26731_ _11681_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_1
X_23943_ _10088_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__buf_4
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35929_ clknet_leaf_475_CLK _04043_ VGND VGND VPWR VPWR registers\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29450_ _13174_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__clkbuf_1
X_26662_ _11644_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ _09550_ registers\[60\]\[17\] _10100_ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__mux2_1
XFILLER_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_805 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_816 _09074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25613_ _11091_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
X_28401_ _12591_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__clkbuf_1
X_29381_ _13137_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_827 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22825_ registers\[60\]\[62\] registers\[61\]\[62\] registers\[62\]\[62\] registers\[63\]\[62\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__mux4_1
X_26593_ _11585_ VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__buf_4
XFILLER_77_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_838 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_849 _09248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28332_ registers\[2\]\[44\] _10397_ _12550_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__mux2_1
X_25544_ _11053_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__clkbuf_1
X_22756_ registers\[32\]\[60\] registers\[33\]\[60\] registers\[34\]\[60\] registers\[35\]\[60\]
+ _07344_ _07345_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__mux4_1
XFILLER_44_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21707_ registers\[12\]\[29\] registers\[13\]\[29\] registers\[14\]\[29\] registers\[15\]\[29\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__mux4_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28263_ registers\[2\]\[11\] _10328_ _12517_ VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__mux2_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25475_ _11017_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_1
X_22687_ registers\[16\]\[57\] registers\[17\]\[57\] registers\[18\]\[57\] registers\[19\]\[57\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__mux4_2
XFILLER_157_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27214_ _11786_ registers\[37\]\[27\] _11958_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__mux2_1
XFILLER_199_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24426_ registers\[57\]\[58\] _10426_ _10410_ VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__mux2_1
X_28194_ _12482_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__clkbuf_1
X_21638_ _08306_ _08309_ _08073_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__o21ba_1
XFILLER_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27145_ _11929_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24357_ net30 VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_382_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_382_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21569_ registers\[24\]\[25\] registers\[25\]\[25\] registers\[26\]\[25\] registers\[27\]\[25\]
+ _08210_ _08211_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__mux4_1
XFILLER_154_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23308_ registers\[9\]\[51\] _09800_ _09798_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__mux2_1
XFILLER_126_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27076_ _11893_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_1
X_24288_ _10333_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26027_ _10747_ registers\[45\]\[8\] _11301_ VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__mux2_1
XFILLER_109_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_134_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23239_ registers\[9\]\[30\] _09753_ _09754_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__mux2_1
XTAP_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1204 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1215 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1226 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17800_ registers\[36\]\[49\] registers\[37\]\[49\] registers\[38\]\[49\] registers\[39\]\[49\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__mux4_1
XANTENNA_1237 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1248 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15992_ registers\[32\]\[0\] registers\[33\]\[0\] registers\[34\]\[0\] registers\[35\]\[0\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _14506_ sky130_fd_sc_hd__mux4_1
XTAP_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_888 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18780_ registers\[24\]\[11\] registers\[25\]\[11\] registers\[26\]\[11\] registers\[27\]\[11\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__mux4_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1259 _00091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27978_ _11738_ registers\[31\]\[4\] _12364_ VGND VGND VPWR VPWR _12369_ sky130_fd_sc_hd__mux2_1
XTAP_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17731_ registers\[56\]\[47\] registers\[57\]\[47\] registers\[58\]\[47\] registers\[59\]\[47\]
+ _04408_ _15885_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__mux4_1
XFILLER_134_1070 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29717_ _13314_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__clkbuf_1
XTAP_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26929_ _11801_ registers\[3\]\[34\] _11793_ VGND VGND VPWR VPWR _11802_ sky130_fd_sc_hd__mux2_1
XFILLER_212_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29648_ registers\[20\]\[61\] _13062_ _13210_ VGND VGND VPWR VPWR _13278_ sky130_fd_sc_hd__mux2_1
X_17662_ registers\[60\]\[45\] registers\[61\]\[45\] registers\[62\]\[45\] registers\[63\]\[45\]
+ _04412_ _15893_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__mux4_1
XFILLER_48_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_1016 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19401_ registers\[52\]\[29\] registers\[53\]\[29\] registers\[54\]\[29\] registers\[55\]\[29\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__mux4_1
X_16613_ registers\[4\]\[15\] registers\[5\]\[15\] registers\[6\]\[15\] registers\[7\]\[15\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _15112_ sky130_fd_sc_hd__mux4_1
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17593_ registers\[56\]\[43\] registers\[57\]\[43\] registers\[58\]\[43\] registers\[59\]\[43\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__mux4_1
XFILLER_169_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29579_ registers\[20\]\[28\] _12993_ _13233_ VGND VGND VPWR VPWR _13242_ sky130_fd_sc_hd__mux2_1
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16544_ _14518_ VGND VGND VPWR VPWR _15045_ sky130_fd_sc_hd__buf_4
X_31610_ registers\[63\]\[30\] net24 _14310_ VGND VGND VPWR VPWR _14311_ sky130_fd_sc_hd__mux2_1
X_19332_ registers\[8\]\[27\] registers\[9\]\[27\] registers\[10\]\[27\] registers\[11\]\[27\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__mux4_1
XFILLER_56_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_962 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32590_ clknet_leaf_72_CLK _00704_ VGND VGND VPWR VPWR registers\[58\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_245_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31541_ _09823_ registers\[6\]\[62\] _14205_ VGND VGND VPWR VPWR _14274_ sky130_fd_sc_hd__mux2_1
X_19263_ registers\[0\]\[25\] registers\[1\]\[25\] registers\[2\]\[25\] registers\[3\]\[25\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__mux4_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16475_ _14796_ _14976_ _14977_ _14799_ VGND VGND VPWR VPWR _14978_ sky130_fd_sc_hd__a22o_1
XFILLER_204_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18214_ _04979_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
X_34260_ clknet_leaf_120_CLK _02374_ VGND VGND VPWR VPWR registers\[32\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31472_ _09751_ registers\[6\]\[29\] _14228_ VGND VGND VPWR VPWR _14238_ sky130_fd_sc_hd__mux2_1
X_19194_ registers\[8\]\[23\] registers\[9\]\[23\] registers\[10\]\[23\] registers\[11\]\[23\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__mux4_1
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33211_ clknet_leaf_299_CLK _01325_ VGND VGND VPWR VPWR registers\[4\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_30423_ _13686_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__clkbuf_1
X_18145_ _04909_ _04912_ _04630_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__o21ba_1
X_34191_ clknet_leaf_132_CLK _02305_ VGND VGND VPWR VPWR registers\[33\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_373_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_373_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18076_ registers\[52\]\[57\] registers\[53\]\[57\] registers\[54\]\[57\] registers\[55\]\[57\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__mux4_1
X_33142_ clknet_leaf_334_CLK _01256_ VGND VGND VPWR VPWR registers\[50\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_30354_ _13650_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17027_ _15198_ _15512_ _15513_ _15204_ VGND VGND VPWR VPWR _15514_ sky130_fd_sc_hd__a22o_1
X_33073_ clknet_leaf_366_CLK _01187_ VGND VGND VPWR VPWR registers\[51\]\[35\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_125_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_125_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30285_ _13613_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__clkbuf_1
X_32024_ clknet_leaf_54_CLK _00202_ VGND VGND VPWR VPWR registers\[62\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18978_ _05720_ _05723_ _05483_ _05484_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__o211a_2
XFILLER_234_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1760 _07379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1771 _10420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ registers\[16\]\[52\] registers\[17\]\[52\] registers\[18\]\[52\] registers\[19\]\[52\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__mux4_1
XANTENNA_1782 _13850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33975_ clknet_leaf_336_CLK _02089_ VGND VGND VPWR VPWR registers\[37\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_239_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35714_ clknet_leaf_241_CLK _03828_ VGND VGND VPWR VPWR registers\[10\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20940_ _07610_ _07617_ _07624_ _07631_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__or4_1
XFILLER_54_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32926_ clknet_leaf_45_CLK _01040_ VGND VGND VPWR VPWR registers\[53\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35645_ clknet_leaf_292_CLK _03759_ VGND VGND VPWR VPWR registers\[11\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20871_ _07564_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
X_32857_ clknet_leaf_66_CLK _00971_ VGND VGND VPWR VPWR registers\[54\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22610_ _09155_ _09252_ _09253_ _09158_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__a22o_1
XFILLER_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31808_ _14414_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23590_ registers\[61\]\[12\] _09683_ _09954_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__mux2_1
X_35576_ clknet_leaf_320_CLK _03690_ VGND VGND VPWR VPWR registers\[12\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_32788_ clknet_leaf_64_CLK _00902_ VGND VGND VPWR VPWR registers\[55\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22541_ _09148_ _09185_ _09186_ _09153_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34527_ clknet_leaf_487_CLK _02641_ VGND VGND VPWR VPWR registers\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31739_ _14378_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25260_ _10800_ registers\[51\]\[33\] _10898_ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__mux2_1
X_22472_ registers\[32\]\[51\] registers\[33\]\[51\] registers\[34\]\[51\] registers\[35\]\[51\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__mux4_1
XFILLER_148_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34458_ clknet_leaf_11_CLK _02572_ VGND VGND VPWR VPWR registers\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_24211_ _09615_ registers\[58\]\[48\] _10277_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__mux2_1
XFILLER_148_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33409_ clknet_leaf_257_CLK _01523_ VGND VGND VPWR VPWR registers\[46\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_21423_ registers\[52\]\[21\] registers\[53\]\[21\] registers\[54\]\[21\] registers\[55\]\[21\]
+ _07919_ _07920_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__mux4_1
X_25191_ _10728_ registers\[51\]\[0\] _10865_ VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_364_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_364_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_34389_ clknet_leaf_97_CLK _02503_ VGND VGND VPWR VPWR registers\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36128_ clknet_leaf_42_CLK _04242_ VGND VGND VPWR VPWR registers\[49\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_24142_ _09546_ registers\[58\]\[15\] _10244_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__mux2_1
XFILLER_136_958 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21354_ registers\[12\]\[19\] registers\[13\]\[19\] registers\[14\]\[19\] registers\[15\]\[19\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__mux4_1
XFILLER_120_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20305_ registers\[40\]\[55\] registers\[41\]\[55\] registers\[42\]\[55\] registers\[43\]\[55\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__mux4_1
XFILLER_200_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_116_CLK clknet_6_20__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_116_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_24073_ _09613_ registers\[5\]\[47\] _10205_ VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__mux2_1
X_36059_ clknet_leaf_35_CLK _04173_ VGND VGND VPWR VPWR registers\[59\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_28950_ registers\[24\]\[17\] _10340_ _12872_ VGND VGND VPWR VPWR _12880_ sky130_fd_sc_hd__mux2_1
XFILLER_100_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21285_ _07963_ _07966_ _07730_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__o21ba_2
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23024_ _09612_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_27901_ _12328_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__clkbuf_1
X_20236_ _06941_ _06946_ _06880_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__o21ba_1
X_28881_ _12843_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_855 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20167_ _05162_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__clkbuf_2
X_27832_ _12291_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__clkbuf_1
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_218_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ _06569_ _06808_ _06811_ _06574_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__a22o_1
X_24975_ _09634_ registers\[53\]\[57\] _10713_ VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__mux2_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27763_ registers\[33\]\[30\] _10367_ _12255_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__mux2_1
XFILLER_218_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29502_ _13201_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__clkbuf_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26714_ _11672_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__clkbuf_1
X_23926_ _10135_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
X_27694_ registers\[34\]\[62\] _10434_ _12150_ VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__mux2_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_602 _05088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_233_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26645_ _11635_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_1
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29433_ _13165_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__clkbuf_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _09533_ registers\[60\]\[9\] _10089_ VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__mux2_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_613 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_624 _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_635 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_646 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22808_ _07343_ _09444_ _09445_ _07353_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__a22o_1
XANTENNA_657 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29364_ _09806_ registers\[22\]\[54\] _13124_ VGND VGND VPWR VPWR _13129_ sky130_fd_sc_hd__mux2_1
X_26576_ _11599_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__clkbuf_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_668 _05396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23788_ _10062_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_232_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_679 _05950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_242_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25527_ _11044_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__clkbuf_1
X_28315_ registers\[2\]\[36\] _10380_ _12539_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__mux2_1
X_22739_ registers\[8\]\[59\] registers\[9\]\[59\] registers\[10\]\[59\] registers\[11\]\[59\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__mux4_1
X_29295_ _09702_ registers\[22\]\[21\] _13091_ VGND VGND VPWR VPWR _13093_ sky130_fd_sc_hd__mux2_1
XFILLER_201_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28246_ registers\[2\]\[3\] _10311_ _12506_ VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__mux2_1
X_16260_ registers\[4\]\[5\] registers\[5\]\[5\] registers\[6\]\[5\] registers\[7\]\[5\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14769_ sky130_fd_sc_hd__mux4_1
XFILLER_125_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25458_ _10862_ registers\[50\]\[63\] _10936_ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__mux2_1
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24409_ _10415_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16191_ _14571_ VGND VGND VPWR VPWR _14702_ sky130_fd_sc_hd__buf_6
X_28177_ _12473_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_355_CLK clknet_6_41__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_355_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25389_ _10936_ VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__buf_4
XFILLER_142_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27128_ _11834_ registers\[38\]\[50\] _11920_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__mux2_1
XFILLER_127_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_107_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_107_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19950_ _06643_ _06652_ _06659_ _06668_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__or4_4
X_27059_ _11884_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18901_ registers\[48\]\[15\] registers\[49\]\[15\] registers\[50\]\[15\] registers\[51\]\[15\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__mux4_1
X_30070_ _13500_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19881_ registers\[20\]\[42\] registers\[21\]\[42\] registers\[22\]\[42\] registers\[23\]\[42\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__mux4_1
XANTENNA_1001 _11828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_214_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1012 _12006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1023 _12505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18832_ _05547_ _05580_ _05581_ _05550_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__a22o_1
XTAP_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1034 _12966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1045 _13281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1056 _13637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1067 _14134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1078 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18763_ registers\[36\]\[11\] registers\[37\]\[11\] registers\[38\]\[11\] registers\[39\]\[11\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__mux4_1
XFILLER_110_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15975_ net67 net68 VGND VGND VPWR VPWR _14489_ sky130_fd_sc_hd__nor2b_4
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1089 _14504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_248_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ registers\[16\]\[46\] registers\[17\]\[46\] registers\[18\]\[46\] registers\[19\]\[46\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__mux4_1
XFILLER_114_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33760_ clknet_leaf_33_CLK _01874_ VGND VGND VPWR VPWR registers\[40\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_30972_ registers\[10\]\[48\] _13035_ _13966_ VGND VGND VPWR VPWR _13975_ sky130_fd_sc_hd__mux2_1
X_18694_ registers\[60\]\[9\] registers\[61\]\[9\] registers\[62\]\[9\] registers\[63\]\[9\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__mux4_1
XFILLER_110_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32711_ clknet_leaf_262_CLK _00825_ VGND VGND VPWR VPWR registers\[57\]\[57\] sky130_fd_sc_hd__dfxtp_1
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17645_ _04289_ _04426_ _04427_ _04292_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__a22o_1
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33691_ clknet_leaf_32_CLK _01805_ VGND VGND VPWR VPWR registers\[41\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35430_ clknet_leaf_461_CLK _03544_ VGND VGND VPWR VPWR registers\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32642_ clknet_leaf_263_CLK _00756_ VGND VGND VPWR VPWR registers\[58\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17576_ registers\[16\]\[42\] registers\[17\]\[42\] registers\[18\]\[42\] registers\[19\]\[42\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__mux4_1
XFILLER_1_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19315_ _06051_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35361_ clknet_leaf_482_CLK _03475_ VGND VGND VPWR VPWR registers\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16527_ registers\[40\]\[13\] registers\[41\]\[13\] registers\[42\]\[13\] registers\[43\]\[13\]
+ _14992_ _14993_ VGND VGND VPWR VPWR _15028_ sky130_fd_sc_hd__mux4_1
X_32573_ clknet_leaf_305_CLK _00687_ VGND VGND VPWR VPWR registers\[5\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34312_ clknet_leaf_245_CLK _02426_ VGND VGND VPWR VPWR registers\[32\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_31524_ _14265_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__clkbuf_1
X_19246_ registers\[40\]\[25\] registers\[41\]\[25\] registers\[42\]\[25\] registers\[43\]\[25\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__mux4_1
X_16458_ _14961_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35292_ clknet_leaf_6_CLK _03406_ VGND VGND VPWR VPWR registers\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34243_ clknet_leaf_250_CLK _02357_ VGND VGND VPWR VPWR registers\[33\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_16389_ _14655_ _14892_ _14893_ _14658_ VGND VGND VPWR VPWR _14894_ sky130_fd_sc_hd__a22o_1
X_31455_ _14229_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19177_ _05912_ _05917_ _05851_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_346_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_346_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18128_ registers\[44\]\[59\] registers\[45\]\[59\] registers\[46\]\[59\] registers\[47\]\[59\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux4_1
X_30406_ _13677_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__clkbuf_1
X_31386_ registers\[7\]\[52\] net48 _14190_ VGND VGND VPWR VPWR _14193_ sky130_fd_sc_hd__mux2_1
X_34174_ clknet_leaf_276_CLK _02288_ VGND VGND VPWR VPWR registers\[34\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_219_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33125_ clknet_leaf_439_CLK _01239_ VGND VGND VPWR VPWR registers\[50\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_18059_ registers\[28\]\[56\] registers\[29\]\[56\] registers\[30\]\[56\] registers\[31\]\[56\]
+ _04706_ _04707_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__mux4_1
X_30337_ _13641_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21070_ registers\[52\]\[11\] registers\[53\]\[11\] registers\[54\]\[11\] registers\[55\]\[11\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__mux4_1
X_30268_ _13604_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__clkbuf_1
X_33056_ clknet_leaf_42_CLK _01170_ VGND VGND VPWR VPWR registers\[51\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20021_ _06737_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__clkbuf_1
X_32007_ clknet_leaf_29_CLK _00180_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
XFILLER_232_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30199_ _13568_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1590 _14518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24760_ _09554_ registers\[54\]\[19\] _10598_ VGND VGND VPWR VPWR _10608_ sky130_fd_sc_hd__mux2_1
XFILLER_67_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21972_ registers\[44\]\[37\] registers\[45\]\[37\] registers\[46\]\[37\] registers\[47\]\[37\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__mux4_1
X_33958_ clknet_leaf_433_CLK _02072_ VGND VGND VPWR VPWR registers\[37\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _09523_ registers\[29\]\[4\] _10017_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__mux2_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32909_ clknet_leaf_140_CLK _01023_ VGND VGND VPWR VPWR registers\[54\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20923_ registers\[52\]\[7\] registers\[53\]\[7\] registers\[54\]\[7\] registers\[55\]\[7\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__mux4_1
XFILLER_227_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24691_ _09622_ registers\[55\]\[51\] _10569_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__mux2_1
XFILLER_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33889_ clknet_leaf_16_CLK _02003_ VGND VGND VPWR VPWR registers\[38\]\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26430_ _10745_ registers\[42\]\[7\] _11514_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__mux2_1
XFILLER_214_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35628_ clknet_leaf_392_CLK _03742_ VGND VGND VPWR VPWR registers\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23642_ registers\[61\]\[37\] _09769_ _09976_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__mux2_1
XFILLER_242_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20854_ _07287_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__buf_6
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_214_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26361_ _11485_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23573_ registers\[61\]\[4\] _09666_ _09943_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__mux2_1
X_35559_ clknet_leaf_460_CLK _03673_ VGND VGND VPWR VPWR registers\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20785_ registers\[52\]\[3\] registers\[53\]\[3\] registers\[54\]\[3\] registers\[55\]\[3\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__mux4_1
X_28100_ _12432_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25312_ _10852_ registers\[51\]\[58\] _10920_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__mux2_1
XFILLER_179_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22524_ registers\[12\]\[52\] registers\[13\]\[52\] registers\[14\]\[52\] registers\[15\]\[52\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__mux4_1
X_29080_ registers\[23\]\[9\] _12953_ _12935_ VGND VGND VPWR VPWR _12954_ sky130_fd_sc_hd__mux2_1
XFILLER_23_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26292_ _11449_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28031_ _12396_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__clkbuf_1
X_25243_ _10783_ registers\[51\]\[25\] _10887_ VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__mux2_1
X_22455_ _07275_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_337_CLK clknet_6_47__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_337_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21406_ _07395_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__clkbuf_4
X_25174_ net55 VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__buf_4
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_194_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22386_ registers\[16\]\[48\] registers\[17\]\[48\] registers\[18\]\[48\] registers\[19\]\[48\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__mux4_1
X_24125_ _09529_ registers\[58\]\[7\] _10233_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__mux2_1
XFILLER_237_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21337_ _07305_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__buf_4
X_29982_ registers\[17\]\[27\] _12991_ _13446_ VGND VGND VPWR VPWR _13454_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28933_ registers\[24\]\[9\] _10323_ _12861_ VGND VGND VPWR VPWR _12871_ sky130_fd_sc_hd__mux2_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24056_ _09596_ registers\[5\]\[39\] _10194_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__mux2_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21268_ _07358_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__buf_4
XFILLER_104_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23007_ net36 VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__clkbuf_4
X_20219_ _06784_ _06928_ _06929_ _06788_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__a22o_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28864_ _11813_ registers\[25\]\[40\] _12834_ VGND VGND VPWR VPWR _12835_ sky130_fd_sc_hd__mux2_1
XFILLER_103_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21199_ _07879_ _07882_ _07711_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__o21ba_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27815_ registers\[33\]\[55\] _10420_ _12277_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__mux2_1
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28795_ _12798_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__clkbuf_1
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24958_ _09617_ registers\[53\]\[49\] _10702_ VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__mux2_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27746_ registers\[33\]\[22\] _10351_ _12244_ VGND VGND VPWR VPWR _12247_ sky130_fd_sc_hd__mux2_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _10126_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
X_27677_ _12210_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_410 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24889_ _09548_ registers\[53\]\[16\] _10669_ VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__mux2_1
XFILLER_209_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_432 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29416_ _13156_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17430_ _15830_ _15902_ _15905_ _15833_ VGND VGND VPWR VPWR _15906_ sky130_fd_sc_hd__a22o_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_443 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26628_ _11626_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_454 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_465 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_476 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29347_ _09788_ registers\[22\]\[46\] _13113_ VGND VGND VPWR VPWR _13120_ sky130_fd_sc_hd__mux2_1
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17361_ registers\[16\]\[36\] registers\[17\]\[36\] registers\[18\]\[36\] registers\[19\]\[36\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _15839_ sky130_fd_sc_hd__mux4_1
XANTENNA_487 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26559_ _11590_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_498 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19100_ _05839_ _05840_ _05841_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a22o_1
X_16312_ _14648_ _14817_ _14818_ _14653_ VGND VGND VPWR VPWR _14819_ sky130_fd_sc_hd__a22o_1
XFILLER_186_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17292_ _15633_ _15770_ _15771_ _15636_ VGND VGND VPWR VPWR _15772_ sky130_fd_sc_hd__a22o_1
XFILLER_202_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29278_ _09685_ registers\[22\]\[13\] _13080_ VGND VGND VPWR VPWR _13084_ sky130_fd_sc_hd__mux2_1
XFILLER_220_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16243_ registers\[44\]\[5\] registers\[45\]\[5\] registers\[46\]\[5\] registers\[47\]\[5\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14752_ sky130_fd_sc_hd__mux4_1
X_19031_ _05501_ _05774_ _05775_ _05506_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__a22o_1
X_28229_ _12500_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_328_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_328_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31240_ registers\[8\]\[47\] net42 _14108_ VGND VGND VPWR VPWR _14116_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16174_ registers\[40\]\[3\] registers\[41\]\[3\] registers\[42\]\[3\] registers\[43\]\[3\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14685_ sky130_fd_sc_hd__mux4_1
XFILLER_220_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput108 net108 VGND VGND VPWR VPWR D1[26] sky130_fd_sc_hd__buf_2
X_31171_ registers\[8\]\[14\] net6 _14075_ VGND VGND VPWR VPWR _14080_ sky130_fd_sc_hd__mux2_1
XFILLER_142_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net119 VGND VGND VPWR VPWR D1[36] sky130_fd_sc_hd__buf_2
XFILLER_141_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30122_ _13527_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19933_ _06647_ _06651_ _06512_ _06513_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__o211a_1
XFILLER_141_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30053_ registers\[17\]\[61\] _13062_ _13423_ VGND VGND VPWR VPWR _13491_ sky130_fd_sc_hd__mux2_1
X_34930_ clknet_leaf_384_CLK _03044_ VGND VGND VPWR VPWR registers\[22\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_19864_ registers\[60\]\[42\] registers\[61\]\[42\] registers\[62\]\[42\] registers\[63\]\[42\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__mux4_1
Xclkbuf_6_2__f_CLK clknet_5_1_0_CLK VGND VGND VPWR VPWR clknet_6_2__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput90 net90 VGND VGND VPWR VPWR D1[0] sky130_fd_sc_hd__buf_2
XFILLER_150_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18815_ _05562_ _05565_ _05494_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__o21ba_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34861_ clknet_leaf_396_CLK _02975_ VGND VGND VPWR VPWR registers\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19795_ registers\[0\]\[40\] registers\[1\]\[40\] registers\[2\]\[40\] registers\[3\]\[40\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__mux4_1
XFILLER_62_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33812_ clknet_leaf_88_CLK _01926_ VGND VGND VPWR VPWR registers\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_18746_ _05146_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__clkbuf_4
XTAP_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34792_ clknet_leaf_452_CLK _02906_ VGND VGND VPWR VPWR registers\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33743_ clknet_leaf_146_CLK _01857_ VGND VGND VPWR VPWR registers\[40\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_18677_ registers\[20\]\[8\] registers\[21\]\[8\] registers\[22\]\[8\] registers\[23\]\[8\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__mux4_1
X_30955_ _13921_ VGND VGND VPWR VPWR _13966_ sky130_fd_sc_hd__buf_4
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17628_ _15884_ _04409_ _04410_ _15890_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a22o_1
XFILLER_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33674_ clknet_leaf_161_CLK _01788_ VGND VGND VPWR VPWR registers\[42\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_30886_ registers\[10\]\[7\] _12949_ _13922_ VGND VGND VPWR VPWR _13930_ sky130_fd_sc_hd__mux2_1
XFILLER_224_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35413_ clknet_leaf_79_CLK _03527_ VGND VGND VPWR VPWR registers\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_32625_ clknet_leaf_367_CLK _00739_ VGND VGND VPWR VPWR registers\[58\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_17559_ _04340_ _04341_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a22o_1
XFILLER_189_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1020 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35344_ clknet_leaf_138_CLK _03458_ VGND VGND VPWR VPWR registers\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20570_ registers\[20\]\[63\] registers\[21\]\[63\] registers\[22\]\[63\] registers\[23\]\[63\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__mux4_1
X_32556_ clknet_leaf_394_CLK _00670_ VGND VGND VPWR VPWR registers\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31507_ _14256_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__clkbuf_1
X_19229_ registers\[0\]\[24\] registers\[1\]\[24\] registers\[2\]\[24\] registers\[3\]\[24\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__mux4_1
X_35275_ clknet_leaf_149_CLK _03389_ VGND VGND VPWR VPWR registers\[17\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_319_CLK clknet_6_39__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_319_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_191_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32487_ clknet_leaf_451_CLK _00601_ VGND VGND VPWR VPWR registers\[60\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22240_ _08891_ _08894_ _08759_ VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__o21ba_1
XFILLER_117_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34226_ clknet_leaf_359_CLK _02340_ VGND VGND VPWR VPWR registers\[33\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31438_ _14220_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34157_ clknet_leaf_321_CLK _02271_ VGND VGND VPWR VPWR registers\[34\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_22171_ registers\[12\]\[42\] registers\[13\]\[42\] registers\[14\]\[42\] registers\[15\]\[42\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__mux4_1
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31369_ registers\[7\]\[44\] net39 _14179_ VGND VGND VPWR VPWR _14184_ sky130_fd_sc_hd__mux2_1
X_33108_ clknet_leaf_70_CLK _01222_ VGND VGND VPWR VPWR registers\[50\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_21122_ registers\[20\]\[12\] registers\[21\]\[12\] registers\[22\]\[12\] registers\[23\]\[12\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__mux4_1
XFILLER_133_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34088_ clknet_leaf_431_CLK _02202_ VGND VGND VPWR VPWR registers\[35\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_801 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33039_ clknet_leaf_75_CLK _01153_ VGND VGND VPWR VPWR registers\[51\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_25930_ _10785_ registers\[46\]\[26\] _11252_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__mux2_1
X_21053_ _07395_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__buf_4
XFILLER_154_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20004_ _06717_ _06718_ _06719_ _06720_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__a22o_1
XFILLER_232_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25861_ _11222_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24812_ _10635_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27600_ registers\[34\]\[17\] _10340_ _12162_ VGND VGND VPWR VPWR _12170_ sky130_fd_sc_hd__mux2_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25792_ _11186_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
X_28580_ _12685_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27531_ _12132_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__clkbuf_1
X_24743_ _10599_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _07366_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__buf_4
XFILLER_243_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20906_ _07386_ _07597_ _07598_ _07396_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__a22o_1
XFILLER_128_1407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27462_ _12096_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__clkbuf_1
X_24674_ _09605_ registers\[55\]\[43\] _10558_ VGND VGND VPWR VPWR _10562_ sky130_fd_sc_hd__mux2_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21886_ _08272_ _08549_ _08550_ _08275_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__a22o_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29201_ registers\[23\]\[48\] _13035_ _13019_ VGND VGND VPWR VPWR _13036_ sky130_fd_sc_hd__mux2_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26413_ _11512_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23625_ registers\[61\]\[29\] _09751_ _09965_ VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__mux2_1
X_20837_ _07528_ _07531_ _07399_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__o21ba_1
X_27393_ registers\[36\]\[48\] _10405_ _12051_ VGND VGND VPWR VPWR _12060_ sky130_fd_sc_hd__mux2_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29132_ net19 VGND VGND VPWR VPWR _12989_ sky130_fd_sc_hd__clkbuf_4
X_26344_ _10793_ registers\[43\]\[30\] _11476_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__mux2_1
X_23556_ _09937_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20768_ registers\[28\]\[2\] registers\[29\]\[2\] registers\[30\]\[2\] registers\[31\]\[2\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__mux4_1
XFILLER_126_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22507_ _09148_ _09151_ _09152_ _09153_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__a22o_1
X_29063_ _12942_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__clkbuf_1
X_26275_ _10860_ registers\[44\]\[62\] _11371_ VGND VGND VPWR VPWR _11440_ sky130_fd_sc_hd__mux2_1
XFILLER_168_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23487_ _09901_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
X_20699_ net76 net75 VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__or2b_4
XFILLER_149_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25226_ _10766_ registers\[51\]\[17\] _10876_ VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__mux2_1
X_28014_ _11774_ registers\[31\]\[21\] _12386_ VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__mux2_1
X_22438_ _09012_ _09085_ _09086_ _09018_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__a22o_1
XFILLER_13_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25157_ _10842_ registers\[52\]\[53\] _10836_ VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__mux2_1
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22369_ _07294_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24108_ _09867_ net83 _09512_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__or3b_1
XFILLER_163_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25088_ net25 VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__buf_4
X_29965_ registers\[17\]\[19\] _12974_ _13435_ VGND VGND VPWR VPWR _13445_ sky130_fd_sc_hd__mux2_1
XFILLER_105_972 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28916_ _12862_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16930_ _15139_ _15418_ _15419_ _15142_ VGND VGND VPWR VPWR _15420_ sky130_fd_sc_hd__a22o_1
X_24039_ _10195_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29896_ registers\[18\]\[50\] _13039_ _13408_ VGND VGND VPWR VPWR _13409_ sky130_fd_sc_hd__mux2_1
XFILLER_132_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28847_ _11797_ registers\[25\]\[32\] _12823_ VGND VGND VPWR VPWR _12826_ sky130_fd_sc_hd__mux2_1
X_16861_ _15349_ _15352_ _15277_ _15278_ VGND VGND VPWR VPWR _15353_ sky130_fd_sc_hd__o211a_1
XFILLER_77_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_889 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18600_ _05141_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__buf_6
XFILLER_19_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19580_ _06304_ _06308_ _06169_ _06170_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__o211a_1
X_28778_ _11584_ _10014_ VGND VGND VPWR VPWR _12789_ sky130_fd_sc_hd__nand2_8
X_16792_ registers\[4\]\[20\] registers\[5\]\[20\] registers\[6\]\[20\] registers\[7\]\[20\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15286_ sky130_fd_sc_hd__mux4_1
XFILLER_237_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18531_ registers\[24\]\[4\] registers\[25\]\[4\] registers\[26\]\[4\] registers\[27\]\[4\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__mux4_1
XFILLER_150_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27729_ registers\[33\]\[14\] _10334_ _12233_ VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__mux2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30740_ _13853_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__clkbuf_1
X_18462_ _05219_ _05222_ _05134_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__o21ba_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_240 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ registers\[48\]\[38\] registers\[49\]\[38\] registers\[50\]\[38\] registers\[51\]\[38\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _15889_ sky130_fd_sc_hd__mux4_1
XANTENNA_273 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18393_ _05092_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__buf_12
X_30671_ registers\[12\]\[33\] _13004_ _13813_ VGND VGND VPWR VPWR _13817_ sky130_fd_sc_hd__mux2_1
XANTENNA_284 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_295 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32410_ clknet_leaf_3_CLK _00524_ VGND VGND VPWR VPWR registers\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ registers\[52\]\[36\] registers\[53\]\[36\] registers\[54\]\[36\] registers\[55\]\[36\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _15822_ sky130_fd_sc_hd__mux4_1
XFILLER_159_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33390_ clknet_leaf_360_CLK _01504_ VGND VGND VPWR VPWR registers\[46\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32341_ clknet_leaf_63_CLK _00455_ VGND VGND VPWR VPWR registers\[61\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17275_ _15541_ _15753_ _15754_ _15547_ VGND VGND VPWR VPWR _15755_ sky130_fd_sc_hd__a22o_1
XFILLER_70_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19014_ _05065_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16226_ registers\[4\]\[4\] registers\[5\]\[4\] registers\[6\]\[4\] registers\[7\]\[4\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14736_ sky130_fd_sc_hd__mux4_1
X_35060_ clknet_leaf_384_CLK _03174_ VGND VGND VPWR VPWR registers\[20\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_32272_ clknet_leaf_113_CLK _00386_ VGND VGND VPWR VPWR registers\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_34011_ clknet_leaf_25_CLK _02125_ VGND VGND VPWR VPWR registers\[36\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_16157_ registers\[0\]\[2\] registers\[1\]\[2\] registers\[2\]\[2\] registers\[3\]\[2\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14669_ sky130_fd_sc_hd__mux4_1
X_31223_ registers\[8\]\[39\] net33 _14097_ VGND VGND VPWR VPWR _14107_ sky130_fd_sc_hd__mux2_1
XFILLER_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16088_ _14592_ VGND VGND VPWR VPWR _14602_ sky130_fd_sc_hd__buf_6
X_31154_ registers\[8\]\[6\] net61 _14064_ VGND VGND VPWR VPWR _14071_ sky130_fd_sc_hd__mux2_1
XFILLER_170_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19916_ _06612_ _06619_ _06628_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__or4_4
X_30105_ registers\[16\]\[21\] _12979_ _13517_ VGND VGND VPWR VPWR _13519_ sky130_fd_sc_hd__mux2_1
XFILLER_64_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35962_ clknet_leaf_304_CLK _04076_ VGND VGND VPWR VPWR registers\[6\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31085_ _14034_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30036_ _13482_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__clkbuf_1
X_34913_ clknet_leaf_489_CLK _03027_ VGND VGND VPWR VPWR registers\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19847_ _06568_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_2
X_35893_ clknet_leaf_323_CLK _04007_ VGND VGND VPWR VPWR registers\[7\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34844_ clknet_leaf_491_CLK _02958_ VGND VGND VPWR VPWR registers\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19778_ registers\[44\]\[40\] registers\[45\]\[40\] registers\[46\]\[40\] registers\[47\]\[40\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__mux4_1
XFILLER_244_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_209_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18729_ _05412_ _05480_ _05481_ _05416_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a22o_1
XFILLER_114_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34775_ clknet_leaf_88_CLK _02889_ VGND VGND VPWR VPWR registers\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1041 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31987_ clknet_leaf_22_CLK _00158_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33726_ clknet_leaf_272_CLK _01840_ VGND VGND VPWR VPWR registers\[41\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_21740_ _07347_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__buf_6
X_30938_ _13957_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33657_ clknet_leaf_339_CLK _01771_ VGND VGND VPWR VPWR registers\[42\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_21671_ registers\[0\]\[28\] registers\[1\]\[28\] registers\[2\]\[28\] registers\[3\]\[28\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__mux4_1
X_30869_ _13920_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_96_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_96_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23410_ _09859_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20622_ registers\[48\]\[0\] registers\[49\]\[0\] registers\[50\]\[0\] registers\[51\]\[0\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__mux4_1
XFILLER_33_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32608_ clknet_leaf_43_CLK _00722_ VGND VGND VPWR VPWR registers\[58\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24390_ _10402_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33588_ clknet_leaf_348_CLK _01702_ VGND VGND VPWR VPWR registers\[43\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23341_ _09822_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
X_35327_ clknet_leaf_196_CLK _03441_ VGND VGND VPWR VPWR registers\[16\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_923 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20553_ registers\[48\]\[63\] registers\[49\]\[63\] registers\[50\]\[63\] registers\[51\]\[63\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__mux4_1
XFILLER_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32539_ clknet_leaf_476_CLK _00653_ VGND VGND VPWR VPWR registers\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26060_ _11327_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__clkbuf_1
X_35258_ clknet_leaf_309_CLK _03372_ VGND VGND VPWR VPWR registers\[17\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_23272_ registers\[9\]\[40\] _09775_ _09776_ VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__mux2_1
X_20484_ _07186_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_138_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25011_ _10743_ registers\[52\]\[6\] _10731_ VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__mux2_1
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22223_ _08812_ _08876_ _08877_ _08815_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__a22o_1
X_34209_ clknet_leaf_43_CLK _02323_ VGND VGND VPWR VPWR registers\[33\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35189_ clknet_leaf_417_CLK _03303_ VGND VGND VPWR VPWR registers\[18\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22154_ _08805_ _08808_ _08809_ _08810_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__a22o_1
XFILLER_238_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21105_ registers\[60\]\[12\] registers\[61\]\[12\] registers\[62\]\[12\] registers\[63\]\[12\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__mux4_1
XFILLER_82_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29750_ registers\[1\]\[45\] _13029_ _13326_ VGND VGND VPWR VPWR _13332_ sky130_fd_sc_hd__mux2_1
XTAP_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26962_ net40 VGND VGND VPWR VPWR _11824_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22085_ _08669_ _08742_ _08743_ _08675_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__a22o_1
XTAP_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_20_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28701_ _11786_ registers\[26\]\[27\] _12741_ VGND VGND VPWR VPWR _12749_ sky130_fd_sc_hd__mux2_1
XFILLER_248_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21036_ registers\[0\]\[10\] registers\[1\]\[10\] registers\[2\]\[10\] registers\[3\]\[10\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__mux4_1
X_25913_ _10768_ registers\[46\]\[18\] _11241_ VGND VGND VPWR VPWR _11250_ sky130_fd_sc_hd__mux2_1
X_29681_ registers\[1\]\[12\] _12960_ _13293_ VGND VGND VPWR VPWR _13296_ sky130_fd_sc_hd__mux2_1
X_26893_ _11777_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_234_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28632_ _12712_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__clkbuf_1
X_25844_ _11213_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28563_ _12676_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__clkbuf_1
X_22987_ _09587_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
X_25775_ _11177_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27514_ _11816_ registers\[35\]\[41\] _12122_ VGND VGND VPWR VPWR _12124_ sky130_fd_sc_hd__mux2_1
X_24726_ _10590_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21938_ registers\[56\]\[36\] registers\[57\]\[36\] registers\[58\]\[36\] registers\[59\]\[36\]
+ _08537_ _08327_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__mux4_1
XFILLER_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28494_ _11849_ registers\[28\]\[57\] _12632_ VGND VGND VPWR VPWR _12640_ sky130_fd_sc_hd__mux2_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27445_ _12087_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24657_ _09588_ registers\[55\]\[35\] _10547_ VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__mux2_1
XFILLER_167_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21869_ registers\[36\]\[34\] registers\[37\]\[34\] registers\[38\]\[34\] registers\[39\]\[34\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_87_CLK clknet_6_18__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_87_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_929 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23608_ _09966_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _09519_ registers\[55\]\[2\] _10514_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__mux2_1
X_27376_ _12006_ VGND VGND VPWR VPWR _12051_ sky130_fd_sc_hd__buf_4
XFILLER_196_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29115_ registers\[23\]\[20\] _12976_ _12977_ VGND VGND VPWR VPWR _12978_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23539_ _09626_ registers\[19\]\[53\] _09925_ VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__mux2_1
XFILLER_169_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26327_ _10777_ registers\[43\]\[22\] _11465_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__mux2_1
XFILLER_11_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17060_ registers\[48\]\[28\] registers\[49\]\[28\] registers\[50\]\[28\] registers\[51\]\[28\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15546_ sky130_fd_sc_hd__mux4_1
X_29046_ registers\[24\]\[63\] _10436_ _12860_ VGND VGND VPWR VPWR _12930_ sky130_fd_sc_hd__mux2_1
X_26258_ _11431_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16011_ _14524_ VGND VGND VPWR VPWR _14525_ sky130_fd_sc_hd__buf_2
XFILLER_195_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25209_ _10749_ registers\[51\]\[9\] _10865_ VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__mux2_1
XFILLER_170_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26189_ _11395_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_15__f_CLK clknet_5_7_0_CLK VGND VGND VPWR VPWR clknet_6_15__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ registers\[24\]\[53\] registers\[25\]\[53\] registers\[26\]\[53\] registers\[27\]\[53\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__mux4_1
XFILLER_139_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29948_ _13436_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_11_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_11_CLK sky130_fd_sc_hd__clkbuf_16
X_19701_ registers\[40\]\[38\] registers\[41\]\[38\] registers\[42\]\[38\] registers\[43\]\[38\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__mux4_1
X_16913_ registers\[32\]\[24\] registers\[33\]\[24\] registers\[34\]\[24\] registers\[35\]\[24\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15403_ sky130_fd_sc_hd__mux4_1
XFILLER_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17893_ registers\[16\]\[51\] registers\[17\]\[51\] registers\[18\]\[51\] registers\[19\]\[51\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__mux4_1
X_29879_ registers\[18\]\[42\] _13023_ _13397_ VGND VGND VPWR VPWR _13400_ sky130_fd_sc_hd__mux2_1
XFILLER_77_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_238_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31910_ _14468_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__clkbuf_1
X_19632_ registers\[32\]\[36\] registers\[33\]\[36\] registers\[34\]\[36\] registers\[35\]\[36\]
+ _06123_ _06124_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__mux4_1
X_16844_ _14496_ VGND VGND VPWR VPWR _15336_ sky130_fd_sc_hd__buf_4
X_32890_ clknet_leaf_287_CLK _01004_ VGND VGND VPWR VPWR registers\[54\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31841_ _14432_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__clkbuf_1
X_19563_ _06269_ _06276_ _06285_ _06292_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__or4_1
XFILLER_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16775_ _14524_ VGND VGND VPWR VPWR _15269_ sky130_fd_sc_hd__buf_2
XFILLER_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18514_ registers\[56\]\[4\] registers\[57\]\[4\] registers\[58\]\[4\] registers\[59\]\[4\]
+ _05272_ _05081_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__mux4_1
X_34560_ clknet_leaf_199_CLK _02674_ VGND VGND VPWR VPWR registers\[28\]\[50\] sky130_fd_sc_hd__dfxtp_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31772_ registers\[59\]\[43\] net38 _14392_ VGND VGND VPWR VPWR _14396_ sky130_fd_sc_hd__mux2_1
X_19494_ _06225_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__buf_2
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33511_ clknet_leaf_60_CLK _01625_ VGND VGND VPWR VPWR registers\[44\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_18445_ registers\[36\]\[2\] registers\[37\]\[2\] registers\[38\]\[2\] registers\[39\]\[2\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__mux4_1
X_30723_ registers\[12\]\[58\] _13056_ _13835_ VGND VGND VPWR VPWR _13844_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34491_ clknet_leaf_301_CLK _02605_ VGND VGND VPWR VPWR registers\[2\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_78_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_78_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36230_ clknet_leaf_121_CLK _00115_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33442_ clknet_leaf_58_CLK _01556_ VGND VGND VPWR VPWR registers\[45\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18376_ _05127_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__buf_4
X_30654_ registers\[12\]\[25\] _12987_ _13802_ VGND VGND VPWR VPWR _13808_ sky130_fd_sc_hd__mux2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_940 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36161_ clknet_leaf_270_CLK _04275_ VGND VGND VPWR VPWR registers\[49\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_17327_ _15638_ _15804_ _15805_ _15643_ VGND VGND VPWR VPWR _15806_ sky130_fd_sc_hd__a22o_1
X_33373_ clknet_leaf_28_CLK _01487_ VGND VGND VPWR VPWR registers\[46\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_30585_ _13771_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35112_ clknet_leaf_458_CLK _03226_ VGND VGND VPWR VPWR registers\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_32324_ clknet_leaf_222_CLK _00438_ VGND VGND VPWR VPWR registers\[19\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_36092_ clknet_leaf_289_CLK _04206_ VGND VGND VPWR VPWR registers\[59\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_17258_ _15633_ _15737_ _15738_ _15636_ VGND VGND VPWR VPWR _15739_ sky130_fd_sc_hd__a22o_1
XFILLER_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16209_ registers\[44\]\[4\] registers\[45\]\[4\] registers\[46\]\[4\] registers\[47\]\[4\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14719_ sky130_fd_sc_hd__mux4_1
X_35043_ clknet_leaf_447_CLK _03157_ VGND VGND VPWR VPWR registers\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_32255_ clknet_leaf_269_CLK _00369_ VGND VGND VPWR VPWR registers\[39\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_17189_ registers\[28\]\[31\] registers\[29\]\[31\] registers\[30\]\[31\] registers\[31\]\[31\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15672_ sky130_fd_sc_hd__mux4_1
XFILLER_143_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31206_ _14098_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32186_ clknet_leaf_466_CLK _00300_ VGND VGND VPWR VPWR registers\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31137_ _14061_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35945_ clknet_leaf_400_CLK _04059_ VGND VGND VPWR VPWR registers\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_31068_ _14025_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22910_ net2 VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__buf_4
XFILLER_96_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30019_ _13473_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35876_ clknet_leaf_467_CLK _03990_ VGND VGND VPWR VPWR registers\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_23890_ _10116_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34827_ clknet_leaf_152_CLK _02941_ VGND VGND VPWR VPWR registers\[24\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_22841_ _07355_ _09476_ _09477_ _07367_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__a22o_1
XFILLER_216_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_225_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25560_ registers\[4\]\[45\] _10399_ _11056_ VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__mux2_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34758_ clknet_leaf_218_CLK _02872_ VGND VGND VPWR VPWR registers\[25\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_22772_ registers\[12\]\[60\] registers\[13\]\[60\] registers\[14\]\[60\] registers\[15\]\[60\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__mux4_1
XFILLER_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24511_ _09580_ registers\[56\]\[31\] _10473_ VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21723_ _07331_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__buf_4
X_33709_ clknet_leaf_330_CLK _01823_ VGND VGND VPWR VPWR registers\[41\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_25491_ registers\[4\]\[12\] _10330_ _11023_ VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__mux2_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34689_ clknet_leaf_222_CLK _02803_ VGND VGND VPWR VPWR registers\[26\]\[51\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_69_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_69_CLK sky130_fd_sc_hd__clkbuf_16
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24442_ _10437_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
X_27230_ _11974_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21654_ _08321_ _08324_ _08054_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__o21ba_1
XFILLER_178_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27161_ _11938_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__clkbuf_1
X_20605_ _07303_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__clkbuf_8
XFILLER_184_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24373_ net36 VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_240_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21585_ registers\[56\]\[26\] registers\[57\]\[26\] registers\[58\]\[26\] registers\[59\]\[26\]
+ _08194_ _07984_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__mux4_1
XFILLER_205_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26112_ _11354_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1088 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23324_ _09811_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
X_20536_ registers\[24\]\[62\] registers\[25\]\[62\] registers\[26\]\[62\] registers\[27\]\[62\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__mux4_1
X_27092_ _11799_ registers\[38\]\[33\] _11898_ VGND VGND VPWR VPWR _11902_ sky130_fd_sc_hd__mux2_1
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26043_ _11318_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23255_ _09765_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20467_ _05149_ _07168_ _07169_ _05159_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__a22o_1
XFILLER_180_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22206_ registers\[4\]\[43\] registers\[5\]\[43\] registers\[6\]\[43\] registers\[7\]\[43\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__mux4_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23186_ _09723_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__clkbuf_1
X_20398_ registers\[44\]\[58\] registers\[45\]\[58\] registers\[46\]\[58\] registers\[47\]\[58\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__mux4_1
Xclkbuf_5_3_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_3_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_106_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29802_ _13359_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__clkbuf_1
XTAP_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22137_ _08615_ _08793_ _08794_ _08618_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__a22o_1
XTAP_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1408 _00177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1419 _00182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput280 net280 VGND VGND VPWR VPWR D3[8] sky130_fd_sc_hd__buf_2
XFILLER_58_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27994_ _12377_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__clkbuf_1
XTAP_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29733_ registers\[1\]\[37\] _13012_ _13315_ VGND VGND VPWR VPWR _13323_ sky130_fd_sc_hd__mux2_1
XTAP_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22068_ registers\[20\]\[39\] registers\[21\]\[39\] registers\[22\]\[39\] registers\[23\]\[39\]
+ _08425_ _08426_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__mux4_1
X_26945_ _11812_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__clkbuf_1
XTAP_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21019_ registers\[44\]\[10\] registers\[45\]\[10\] registers\[46\]\[10\] registers\[47\]\[10\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__mux4_1
X_29664_ registers\[1\]\[4\] _12943_ _13282_ VGND VGND VPWR VPWR _13287_ sky130_fd_sc_hd__mux2_1
XTAP_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26876_ _11765_ registers\[3\]\[17\] _11751_ VGND VGND VPWR VPWR _11766_ sky130_fd_sc_hd__mux2_1
XFILLER_102_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28615_ _11834_ registers\[27\]\[50\] _12703_ VGND VGND VPWR VPWR _12704_ sky130_fd_sc_hd__mux2_1
X_25827_ _10817_ registers\[47\]\[41\] _11203_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__mux2_1
X_29595_ _13250_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28546_ _12667_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__clkbuf_1
X_16560_ registers\[32\]\[14\] registers\[33\]\[14\] registers\[34\]\[14\] registers\[35\]\[14\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _15060_ sky130_fd_sc_hd__mux4_1
X_25758_ _11168_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24709_ _09640_ registers\[55\]\[60\] _10513_ VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__mux2_1
XFILLER_203_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28477_ _11832_ registers\[28\]\[49\] _12621_ VGND VGND VPWR VPWR _12631_ sky130_fd_sc_hd__mux2_1
XFILLER_16_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16491_ _14496_ VGND VGND VPWR VPWR _14993_ sky130_fd_sc_hd__buf_4
X_25689_ _11131_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18230_ registers\[0\]\[62\] registers\[1\]\[62\] registers\[2\]\[62\] registers\[3\]\[62\]
+ _14621_ _14622_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__mux4_1
XFILLER_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27428_ _11728_ registers\[35\]\[0\] _12078_ VGND VGND VPWR VPWR _12079_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_0_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18161_ _04924_ _04927_ _14524_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__o21ba_1
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27359_ _12042_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17112_ registers\[16\]\[29\] registers\[17\]\[29\] registers\[18\]\[29\] registers\[19\]\[29\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15597_ sky130_fd_sc_hd__mux4_1
X_18092_ _04858_ _04861_ _04644_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__o21ba_1
X_30370_ _13658_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29029_ _12921_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__clkbuf_1
X_17043_ registers\[20\]\[27\] registers\[21\]\[27\] registers\[22\]\[27\] registers\[23\]\[27\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15530_ sky130_fd_sc_hd__mux4_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32040_ clknet_leaf_436_CLK _00218_ VGND VGND VPWR VPWR registers\[62\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1084 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_1054 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18994_ _05739_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17945_ _04715_ _04718_ _04611_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__o21ba_1
XFILLER_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33991_ clknet_leaf_236_CLK _02105_ VGND VGND VPWR VPWR registers\[37\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_239_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35730_ clknet_leaf_106_CLK _03844_ VGND VGND VPWR VPWR registers\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_32942_ clknet_leaf_368_CLK _01056_ VGND VGND VPWR VPWR registers\[53\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17876_ _04340_ _04650_ _04651_ _04343_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a22o_1
XFILLER_241_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19615_ registers\[8\]\[35\] registers\[9\]\[35\] registers\[10\]\[35\] registers\[11\]\[35\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__mux4_1
X_35661_ clknet_leaf_146_CLK _03775_ VGND VGND VPWR VPWR registers\[11\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16827_ registers\[0\]\[21\] registers\[1\]\[21\] registers\[2\]\[21\] registers\[3\]\[21\]
+ _15281_ _15282_ VGND VGND VPWR VPWR _15320_ sky130_fd_sc_hd__mux4_1
X_32873_ clknet_leaf_423_CLK _00987_ VGND VGND VPWR VPWR registers\[54\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_242_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34612_ clknet_leaf_413_CLK _02726_ VGND VGND VPWR VPWR registers\[27\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_207_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31824_ _14423_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__clkbuf_1
X_19546_ _06272_ _06275_ _06169_ _06170_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__o211a_1
X_35592_ clknet_leaf_156_CLK _03706_ VGND VGND VPWR VPWR registers\[12\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_16758_ registers\[24\]\[19\] registers\[25\]\[19\] registers\[26\]\[19\] registers\[27\]\[19\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15253_ sky130_fd_sc_hd__mux4_1
XFILLER_207_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34543_ clknet_leaf_395_CLK _02657_ VGND VGND VPWR VPWR registers\[28\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_206_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31755_ registers\[59\]\[35\] net29 _14381_ VGND VGND VPWR VPWR _14387_ sky130_fd_sc_hd__mux2_1
X_19477_ _06098_ _06207_ _06208_ _06102_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__a22o_1
XFILLER_59_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16689_ registers\[28\]\[17\] registers\[29\]\[17\] registers\[30\]\[17\] registers\[31\]\[17\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15186_ sky130_fd_sc_hd__mux4_1
XFILLER_59_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_895 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30706_ _13779_ VGND VGND VPWR VPWR _13835_ sky130_fd_sc_hd__buf_4
X_18428_ registers\[16\]\[1\] registers\[17\]\[1\] registers\[18\]\[1\] registers\[19\]\[1\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux4_1
X_34474_ clknet_leaf_458_CLK _02588_ VGND VGND VPWR VPWR registers\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_31686_ registers\[59\]\[2\] net23 _14348_ VGND VGND VPWR VPWR _14351_ sky130_fd_sc_hd__mux2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36213_ clknet_leaf_115_CLK _00096_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dfxtp_1
XFILLER_148_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33425_ clknet_leaf_130_CLK _01539_ VGND VGND VPWR VPWR registers\[45\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_18359_ _05044_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__buf_12
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30637_ registers\[12\]\[17\] _12970_ _13791_ VGND VGND VPWR VPWR _13799_ sky130_fd_sc_hd__mux2_1
XFILLER_30_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36144_ clknet_leaf_365_CLK _04258_ VGND VGND VPWR VPWR registers\[49\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_33356_ clknet_leaf_176_CLK _01470_ VGND VGND VPWR VPWR registers\[47\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_21370_ _07331_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__buf_4
XFILLER_108_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30568_ _13762_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20321_ _06717_ _07027_ _07028_ _06720_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__a22o_1
X_32307_ clknet_leaf_409_CLK _00421_ VGND VGND VPWR VPWR registers\[19\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36075_ clknet_leaf_420_CLK _04189_ VGND VGND VPWR VPWR registers\[59\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_33287_ clknet_leaf_260_CLK _01401_ VGND VGND VPWR VPWR registers\[48\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_30499_ _13726_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23040_ _09623_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
X_35026_ clknet_leaf_101_CLK _03140_ VGND VGND VPWR VPWR registers\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_20252_ _06958_ _06961_ _06855_ _06856_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__o211a_1
X_32238_ clknet_leaf_357_CLK _00352_ VGND VGND VPWR VPWR registers\[39\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20183_ _06784_ _06893_ _06894_ _06788_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__a22o_1
X_32169_ clknet_leaf_79_CLK _00283_ VGND VGND VPWR VPWR registers\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_61__f_CLK clknet_5_30_0_CLK VGND VGND VPWR VPWR clknet_6_61__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_24991_ _10512_ _10729_ VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__nand2_8
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26730_ registers\[40\]\[20\] _10346_ _11680_ VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__mux2_1
XFILLER_229_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23942_ _10143_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35928_ clknet_leaf_474_CLK _04042_ VGND VGND VPWR VPWR registers\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26661_ _10840_ registers\[41\]\[52\] _11641_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__mux2_1
X_23873_ _10107_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35859_ clknet_leaf_78_CLK _03973_ VGND VGND VPWR VPWR registers\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28400_ _11755_ registers\[28\]\[12\] _12588_ VGND VGND VPWR VPWR _12591_ sky130_fd_sc_hd__mux2_1
XFILLER_38_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22824_ _07372_ _09459_ _09460_ _07382_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__a22o_1
XANTENNA_806 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25612_ registers\[48\]\[4\] _10313_ _11086_ VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__mux2_1
XANTENNA_817 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29380_ _09823_ registers\[22\]\[62\] _13068_ VGND VGND VPWR VPWR _13137_ sky130_fd_sc_hd__mux2_1
XANTENNA_828 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26592_ _11607_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_839 _09184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28331_ _12554_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22755_ registers\[40\]\[60\] registers\[41\]\[60\] registers\[42\]\[60\] registers\[43\]\[60\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__mux4_1
X_25543_ registers\[4\]\[37\] _10382_ _11045_ VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__mux2_1
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_213_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21706_ _08267_ _08374_ _08375_ _08270_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__a22o_1
XFILLER_198_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25474_ registers\[4\]\[4\] _10313_ _11012_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__mux2_1
X_28262_ _12518_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__clkbuf_1
X_22686_ registers\[24\]\[57\] registers\[25\]\[57\] registers\[26\]\[57\] registers\[27\]\[57\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__mux4_1
XFILLER_212_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24425_ net54 VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__buf_4
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27213_ _11965_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21637_ _08272_ _08307_ _08308_ _08275_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__a22o_1
XFILLER_90_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28193_ _11818_ registers\[30\]\[42\] _12479_ VGND VGND VPWR VPWR _12482_ sky130_fd_sc_hd__mux2_1
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27144_ _11851_ registers\[38\]\[58\] _11920_ VGND VGND VPWR VPWR _11929_ sky130_fd_sc_hd__mux2_1
XFILLER_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24356_ _10379_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
X_21568_ _08238_ _08241_ _08073_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__o21ba_1
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23307_ net47 VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__buf_4
XFILLER_165_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20519_ registers\[36\]\[62\] registers\[37\]\[62\] registers\[38\]\[62\] registers\[39\]\[62\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__mux4_1
XFILLER_153_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27075_ _11782_ registers\[38\]\[25\] _11887_ VGND VGND VPWR VPWR _11893_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24287_ registers\[57\]\[13\] _10332_ _10326_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__mux2_1
X_21499_ registers\[12\]\[23\] registers\[13\]\[23\] registers\[14\]\[23\] registers\[15\]\[23\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__mux4_1
XFILLER_181_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26026_ _11309_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23238_ _09708_ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__buf_4
XFILLER_5_969 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23169_ registers\[9\]\[4\] _09666_ _09709_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__mux2_1
XANTENNA_1205 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1216 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1227 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1238 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15991_ _14504_ VGND VGND VPWR VPWR _14505_ sky130_fd_sc_hd__buf_4
XTAP_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27977_ _12368_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1249 _00090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _04504_ _04509_ _15955_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__o21ba_1
X_29716_ registers\[1\]\[29\] _12995_ _13304_ VGND VGND VPWR VPWR _13314_ sky130_fd_sc_hd__mux2_1
XFILLER_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26928_ net28 VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__clkbuf_4
XTAP_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29647_ _13277_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__clkbuf_1
XTAP_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _15884_ _04441_ _04442_ _15890_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__a22o_1
XFILLER_236_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26859_ _11754_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19400_ registers\[60\]\[29\] registers\[61\]\[29\] registers\[62\]\[29\] registers\[63\]\[29\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16612_ registers\[12\]\[15\] registers\[13\]\[15\] registers\[14\]\[15\] registers\[15\]\[15\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15111_ sky130_fd_sc_hd__mux4_1
X_17592_ _04372_ _04375_ _15955_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__o21ba_1
X_29578_ _13241_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19331_ _06063_ _06066_ _05826_ _05827_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o211a_1
XFILLER_189_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28529_ _12658_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__clkbuf_1
X_16543_ _14796_ _15042_ _15043_ _14799_ VGND VGND VPWR VPWR _15044_ sky130_fd_sc_hd__a22o_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_232_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31540_ _14273_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_206_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19262_ registers\[8\]\[25\] registers\[9\]\[25\] registers\[10\]\[25\] registers\[11\]\[25\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__mux4_1
X_16474_ registers\[0\]\[11\] registers\[1\]\[11\] registers\[2\]\[11\] registers\[3\]\[11\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _14977_ sky130_fd_sc_hd__mux4_1
X_18213_ _04957_ _04964_ _04971_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__or4_4
X_31471_ _14237_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19193_ _05929_ _05932_ _05826_ _05827_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__o211a_1
XFILLER_129_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33210_ clknet_leaf_304_CLK _01324_ VGND VGND VPWR VPWR registers\[4\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_18144_ _14511_ _04910_ _04911_ _14517_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__a22o_1
XFILLER_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30422_ _09782_ registers\[14\]\[43\] _13682_ VGND VGND VPWR VPWR _13686_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34190_ clknet_leaf_131_CLK _02304_ VGND VGND VPWR VPWR registers\[33\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_1146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33141_ clknet_leaf_328_CLK _01255_ VGND VGND VPWR VPWR registers\[50\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_18075_ registers\[60\]\[57\] registers\[61\]\[57\] registers\[62\]\[57\] registers\[63\]\[57\]
+ _04755_ _04549_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__mux4_1
X_30353_ _09678_ registers\[14\]\[10\] _13649_ VGND VGND VPWR VPWR _13650_ sky130_fd_sc_hd__mux2_1
XFILLER_32_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17026_ registers\[48\]\[27\] registers\[49\]\[27\] registers\[50\]\[27\] registers\[51\]\[27\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15513_ sky130_fd_sc_hd__mux4_1
XFILLER_109_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33072_ clknet_leaf_366_CLK _01186_ VGND VGND VPWR VPWR registers\[51\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30284_ registers\[15\]\[42\] _13023_ _13610_ VGND VGND VPWR VPWR _13613_ sky130_fd_sc_hd__mux2_1
XFILLER_217_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32023_ clknet_leaf_62_CLK _00201_ VGND VGND VPWR VPWR registers\[62\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _05412_ _05721_ _05722_ _05416_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__a22o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1750 _06309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1761 _07379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17928_ registers\[24\]\[52\] registers\[25\]\[52\] registers\[26\]\[52\] registers\[27\]\[52\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux4_1
XFILLER_234_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_932 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1772 _11300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33974_ clknet_leaf_336_CLK _02088_ VGND VGND VPWR VPWR registers\[37\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1783 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35713_ clknet_leaf_240_CLK _03827_ VGND VGND VPWR VPWR registers\[10\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32925_ clknet_leaf_54_CLK _01039_ VGND VGND VPWR VPWR registers\[53\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17859_ _04632_ _04633_ _04634_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__a22o_1
XFILLER_67_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20870_ _07540_ _07547_ _07556_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__or4_2
X_35644_ clknet_leaf_300_CLK _03758_ VGND VGND VPWR VPWR registers\[11\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_32856_ clknet_leaf_52_CLK _00970_ VGND VGND VPWR VPWR registers\[54\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31807_ registers\[59\]\[60\] net57 _14347_ VGND VGND VPWR VPWR _14414_ sky130_fd_sc_hd__mux2_1
X_19529_ _06187_ _06258_ _06259_ _06192_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__a22o_1
XFILLER_228_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35575_ clknet_leaf_319_CLK _03689_ VGND VGND VPWR VPWR registers\[12\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32787_ clknet_leaf_182_CLK _00901_ VGND VGND VPWR VPWR registers\[55\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22540_ registers\[32\]\[53\] registers\[33\]\[53\] registers\[34\]\[53\] registers\[35\]\[53\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__mux4_1
X_34526_ clknet_leaf_490_CLK _02640_ VGND VGND VPWR VPWR registers\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31738_ registers\[59\]\[27\] net20 _14370_ VGND VGND VPWR VPWR _14378_ sky130_fd_sc_hd__mux2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22471_ registers\[40\]\[51\] registers\[41\]\[51\] registers\[42\]\[51\] registers\[43\]\[51\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__mux4_1
X_34457_ clknet_leaf_11_CLK _02571_ VGND VGND VPWR VPWR registers\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31669_ _14341_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24210_ _10285_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
X_33408_ clknet_leaf_257_CLK _01522_ VGND VGND VPWR VPWR registers\[46\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21422_ registers\[60\]\[21\] registers\[61\]\[21\] registers\[62\]\[21\] registers\[63\]\[21\]
+ _07855_ _07992_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__mux4_1
XFILLER_182_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25190_ _10864_ VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__clkbuf_4
X_34388_ clknet_leaf_94_CLK _02502_ VGND VGND VPWR VPWR registers\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36127_ clknet_leaf_38_CLK _04241_ VGND VGND VPWR VPWR registers\[49\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_24141_ _10249_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__clkbuf_1
X_33339_ clknet_leaf_278_CLK _01453_ VGND VGND VPWR VPWR registers\[47\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_21353_ _07924_ _08031_ _08032_ _07927_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__a22o_1
XFILLER_194_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20304_ _07012_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__buf_4
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24072_ _10212_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_36058_ clknet_leaf_83_CLK _04172_ VGND VGND VPWR VPWR registers\[59\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_21284_ _07929_ _07964_ _07965_ _07932_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__a22o_1
XFILLER_190_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35009_ clknet_leaf_202_CLK _03123_ VGND VGND VPWR VPWR registers\[21\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_23023_ _09611_ registers\[62\]\[46\] _09599_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__mux2_1
XFILLER_144_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27900_ registers\[32\]\[31\] _10370_ _12326_ VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__mux2_1
X_20235_ _06873_ _06944_ _06945_ _06878_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__a22o_1
X_28880_ _11830_ registers\[25\]\[48\] _12834_ VGND VGND VPWR VPWR _12843_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27831_ registers\[33\]\[63\] _10436_ _12221_ VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__mux2_1
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _06873_ _06874_ _06877_ _06878_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__a22o_1
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27762_ _12221_ VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__buf_4
X_20097_ registers\[32\]\[49\] registers\[33\]\[49\] registers\[34\]\[49\] registers\[35\]\[49\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__mux4_1
X_24974_ _10720_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29501_ _09808_ registers\[21\]\[55\] _13195_ VGND VGND VPWR VPWR _13201_ sky130_fd_sc_hd__mux2_1
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26713_ registers\[40\]\[12\] _10330_ _11669_ VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__mux2_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23925_ _09601_ registers\[60\]\[41\] _10133_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__mux2_1
XFILLER_218_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27693_ _12218_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29432_ _09717_ registers\[21\]\[22\] _13162_ VGND VGND VPWR VPWR _13165_ sky130_fd_sc_hd__mux2_1
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_603 _05095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26644_ _10823_ registers\[41\]\[44\] _11630_ VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__mux2_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23856_ _10098_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_614 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_625 _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_636 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22807_ registers\[16\]\[61\] registers\[17\]\[61\] registers\[18\]\[61\] registers\[19\]\[61\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__mux4_1
X_29363_ _13128_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_647 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26575_ _10754_ registers\[41\]\[11\] _11597_ VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__mux2_1
XANTENNA_658 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ registers\[0\]\[9\] registers\[1\]\[9\] registers\[2\]\[9\] registers\[3\]\[9\]
+ _07348_ _07350_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__mux4_1
XANTENNA_669 _05396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23787_ _09598_ registers\[29\]\[40\] _10061_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__mux2_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28314_ _12545_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25526_ registers\[4\]\[29\] _10365_ _11034_ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__mux2_1
X_22738_ _09374_ _09377_ _09091_ _09092_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__o211a_1
X_29294_ _13092_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1067 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28245_ _12509_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22669_ registers\[36\]\[57\] registers\[37\]\[57\] registers\[38\]\[57\] registers\[39\]\[57\]
+ _07357_ _07359_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__mux4_1
XFILLER_199_1105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25457_ _11005_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24408_ registers\[57\]\[52\] _10414_ _10410_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__mux2_1
XFILLER_138_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16190_ _14558_ _14699_ _14700_ _14568_ VGND VGND VPWR VPWR _14701_ sky130_fd_sc_hd__a22o_1
X_28176_ _11801_ registers\[30\]\[34\] _12468_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__mux2_1
XFILLER_154_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25388_ _10969_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27127_ _11864_ VGND VGND VPWR VPWR _11920_ sky130_fd_sc_hd__buf_4
XFILLER_103_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24339_ _10304_ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__clkbuf_8
XFILLER_193_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27058_ _11765_ registers\[38\]\[17\] _11876_ VGND VGND VPWR VPWR _11884_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18900_ registers\[56\]\[15\] registers\[57\]\[15\] registers\[58\]\[15\] registers\[59\]\[15\]
+ _05615_ _05405_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__mux4_1
X_26009_ _10015_ _11157_ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__nand2_8
X_19880_ registers\[28\]\[42\] registers\[29\]\[42\] registers\[30\]\[42\] registers\[31\]\[42\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__mux4_1
XFILLER_84_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1002 _11830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18831_ registers\[36\]\[13\] registers\[37\]\[13\] registers\[38\]\[13\] registers\[39\]\[13\]
+ _05370_ _05371_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__mux4_1
XANTENNA_1013 _12077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1024 _12505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1035 _13012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1046 _13281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1057 _13779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18762_ registers\[44\]\[11\] registers\[45\]\[11\] registers\[46\]\[11\] registers\[47\]\[11\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__mux4_1
XANTENNA_1068 _14205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1079 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _14532_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__buf_4
XTAP_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30971_ _13974_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__clkbuf_1
X_18693_ _05404_ _05445_ _05446_ _05410_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a22o_1
XFILLER_64_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32710_ clknet_leaf_262_CLK _00824_ VGND VGND VPWR VPWR registers\[57\]\[56\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_291_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_291_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ registers\[16\]\[44\] registers\[17\]\[44\] registers\[18\]\[44\] registers\[19\]\[44\]
+ _15837_ _15838_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__mux4_1
XFILLER_236_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33690_ clknet_leaf_32_CLK _01804_ VGND VGND VPWR VPWR registers\[41\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32641_ clknet_leaf_266_CLK _00755_ VGND VGND VPWR VPWR registers\[58\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17575_ registers\[24\]\[42\] registers\[25\]\[42\] registers\[26\]\[42\] registers\[27\]\[42\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__mux4_1
X_19314_ _06021_ _06030_ _06041_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__or4_4
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35360_ clknet_leaf_482_CLK _03474_ VGND VGND VPWR VPWR registers\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16526_ _15027_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32572_ clknet_leaf_299_CLK _00686_ VGND VGND VPWR VPWR registers\[5\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34311_ clknet_leaf_244_CLK _02425_ VGND VGND VPWR VPWR registers\[32\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31523_ _09804_ registers\[6\]\[53\] _14261_ VGND VGND VPWR VPWR _14265_ sky130_fd_sc_hd__mux2_1
X_19245_ _05983_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__clkbuf_1
X_35291_ clknet_leaf_6_CLK _03405_ VGND VGND VPWR VPWR registers\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_16457_ _14927_ _14936_ _14946_ _14960_ VGND VGND VPWR VPWR _14961_ sky130_fd_sc_hd__or4_2
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34242_ clknet_leaf_249_CLK _02356_ VGND VGND VPWR VPWR registers\[33\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_31454_ _09699_ registers\[6\]\[20\] _14228_ VGND VGND VPWR VPWR _14229_ sky130_fd_sc_hd__mux2_1
X_19176_ _05844_ _05915_ _05916_ _05849_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__a22o_1
X_16388_ registers\[36\]\[9\] registers\[37\]\[9\] registers\[38\]\[9\] registers\[39\]\[9\]
+ _14821_ _14822_ VGND VGND VPWR VPWR _14893_ sky130_fd_sc_hd__mux4_1
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18127_ _04676_ _04893_ _04894_ _04681_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__a22o_1
X_30405_ _09764_ registers\[14\]\[35\] _13671_ VGND VGND VPWR VPWR _13677_ sky130_fd_sc_hd__mux2_1
X_34173_ clknet_leaf_276_CLK _02287_ VGND VGND VPWR VPWR registers\[34\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_31385_ _14192_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33124_ clknet_leaf_440_CLK _01238_ VGND VGND VPWR VPWR registers\[50\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_18058_ _04632_ _04827_ _04828_ _04635_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__a22o_1
X_30336_ _09662_ registers\[14\]\[2\] _13638_ VGND VGND VPWR VPWR _13641_ sky130_fd_sc_hd__mux2_1
XFILLER_172_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17009_ _15290_ _15493_ _15496_ _15293_ VGND VGND VPWR VPWR _15497_ sky130_fd_sc_hd__a22o_1
XFILLER_119_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33055_ clknet_leaf_36_CLK _01169_ VGND VGND VPWR VPWR registers\[51\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_30267_ registers\[15\]\[34\] _13006_ _13599_ VGND VGND VPWR VPWR _13604_ sky130_fd_sc_hd__mux2_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20020_ _06707_ _06716_ _06727_ _06736_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__or4_4
X_32006_ clknet_leaf_28_CLK _00179_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30198_ registers\[15\]\[1\] _12937_ _13566_ VGND VGND VPWR VPWR _13568_ sky130_fd_sc_hd__mux2_1
XFILLER_80_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_230_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1580 _13921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1591 _14539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21971_ _08462_ _08631_ _08632_ _08467_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__a22o_1
X_33957_ clknet_leaf_433_CLK _02071_ VGND VGND VPWR VPWR registers\[37\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_282_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_282_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23710_ _10021_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
X_20922_ registers\[60\]\[7\] registers\[61\]\[7\] registers\[62\]\[7\] registers\[63\]\[7\]
+ _07512_ _07329_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__mux4_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32908_ clknet_leaf_142_CLK _01022_ VGND VGND VPWR VPWR registers\[54\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_24690_ _10570_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33888_ clknet_leaf_16_CLK _02002_ VGND VGND VPWR VPWR registers\[38\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32839_ clknet_leaf_196_CLK _00953_ VGND VGND VPWR VPWR registers\[55\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_20853_ _07543_ _07546_ _07339_ _07341_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__o211a_1
X_35627_ clknet_leaf_399_CLK _03741_ VGND VGND VPWR VPWR registers\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _09983_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_214_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23572_ _09947_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
X_26360_ _10810_ registers\[43\]\[38\] _11476_ VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__mux2_1
X_20784_ registers\[60\]\[3\] registers\[61\]\[3\] registers\[62\]\[3\] registers\[63\]\[3\]
+ _07327_ _07329_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__mux4_1
X_35558_ clknet_leaf_461_CLK _03672_ VGND VGND VPWR VPWR registers\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22523_ _08953_ _09168_ _09169_ _08956_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__a22o_1
XFILLER_210_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25311_ _10928_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__clkbuf_1
X_34509_ clknet_leaf_147_CLK _02623_ VGND VGND VPWR VPWR registers\[2\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_26291_ _10741_ registers\[43\]\[5\] _11443_ VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__mux2_1
XFILLER_194_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35489_ clknet_leaf_483_CLK _03603_ VGND VGND VPWR VPWR registers\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28030_ _11790_ registers\[31\]\[29\] _12386_ VGND VGND VPWR VPWR _12396_ sky130_fd_sc_hd__mux2_1
X_22454_ _09098_ _09101_ _09102_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__o21ba_1
X_25242_ _10892_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_926 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21405_ registers\[20\]\[20\] registers\[21\]\[20\] registers\[22\]\[20\] registers\[23\]\[20\]
+ _08082_ _08083_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__mux4_1
X_25173_ _10853_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__clkbuf_1
X_22385_ registers\[24\]\[48\] registers\[25\]\[48\] registers\[26\]\[48\] registers\[27\]\[48\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__mux4_1
XFILLER_136_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24124_ _10240_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21336_ _07303_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__buf_4
XFILLER_194_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29981_ _13453_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1046 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_237_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28932_ _12870_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__clkbuf_1
X_24055_ _10203_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
X_21267_ _07356_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__buf_4
XFILLER_235_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23006_ _09600_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
X_20218_ registers\[52\]\[52\] registers\[53\]\[52\] registers\[54\]\[52\] registers\[55\]\[52\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__mux4_1
X_28863_ _12789_ VGND VGND VPWR VPWR _12834_ sky130_fd_sc_hd__clkbuf_8
XFILLER_132_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21198_ _07783_ _07880_ _07881_ _07786_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__a22o_1
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27814_ _12282_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__clkbuf_1
X_20149_ _06717_ _06858_ _06861_ _06720_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__a22o_1
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28794_ _11744_ registers\[25\]\[7\] _12790_ VGND VGND VPWR VPWR _12798_ sky130_fd_sc_hd__mux2_1
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27745_ _12246_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_218_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24957_ _10711_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__clkbuf_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_273_CLK clknet_6_59__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_273_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23908_ _09584_ registers\[60\]\[33\] _10122_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__mux2_1
XFILLER_46_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27676_ registers\[34\]\[53\] _10416_ _12206_ VGND VGND VPWR VPWR _12210_ sky130_fd_sc_hd__mux2_1
XFILLER_131_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24888_ _10675_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__clkbuf_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29415_ _09687_ registers\[21\]\[14\] _13151_ VGND VGND VPWR VPWR _13156_ sky130_fd_sc_hd__mux2_1
XFILLER_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_433 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26627_ _10806_ registers\[41\]\[36\] _11619_ VGND VGND VPWR VPWR _11626_ sky130_fd_sc_hd__mux2_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23839_ _09510_ registers\[60\]\[0\] _10089_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__mux2_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_444 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_455 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_466 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _14532_ VGND VGND VPWR VPWR _15838_ sky130_fd_sc_hd__buf_4
X_29346_ _13119_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_477 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26558_ _10737_ registers\[41\]\[3\] _11586_ VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__mux2_1
XFILLER_25_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_488 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_499 _00167_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16311_ registers\[32\]\[7\] registers\[33\]\[7\] registers\[34\]\[7\] registers\[35\]\[7\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14818_ sky130_fd_sc_hd__mux4_1
XFILLER_213_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_876 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25509_ _11035_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29277_ _13083_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__clkbuf_1
X_17291_ registers\[16\]\[34\] registers\[17\]\[34\] registers\[18\]\[34\] registers\[19\]\[34\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15771_ sky130_fd_sc_hd__mux4_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26489_ _10804_ registers\[42\]\[35\] _11547_ VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__mux2_1
XFILLER_207_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_1470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_202_988 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19030_ registers\[20\]\[18\] registers\[21\]\[18\] registers\[22\]\[18\] registers\[23\]\[18\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__mux4_1
X_16242_ _14648_ _14749_ _14750_ _14653_ VGND VGND VPWR VPWR _14751_ sky130_fd_sc_hd__a22o_1
X_28228_ _11853_ registers\[30\]\[59\] _12490_ VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__mux2_1
XFILLER_185_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16173_ _14684_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28159_ _11784_ registers\[30\]\[26\] _12457_ VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__mux2_1
XFILLER_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR D1[27] sky130_fd_sc_hd__buf_2
X_31170_ _14079_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30121_ registers\[16\]\[29\] _12995_ _13517_ VGND VGND VPWR VPWR _13527_ sky130_fd_sc_hd__mux2_1
XFILLER_99_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19932_ _06441_ _06649_ _06650_ _06445_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__a22o_1
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30052_ _13490_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__clkbuf_1
X_19863_ _06433_ _06582_ _06583_ _06439_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__a22o_1
XFILLER_95_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput91 net91 VGND VGND VPWR VPWR D1[10] sky130_fd_sc_hd__buf_2
XFILLER_214_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_214_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18814_ _05350_ _05563_ _05564_ _05353_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a22o_1
XTAP_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19794_ _05122_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34860_ clknet_leaf_395_CLK _02974_ VGND VGND VPWR VPWR registers\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_237_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33811_ clknet_leaf_105_CLK _01925_ VGND VGND VPWR VPWR registers\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_18745_ registers\[16\]\[10\] registers\[17\]\[10\] registers\[18\]\[10\] registers\[19\]\[10\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__mux4_1
XFILLER_62_1182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34791_ clknet_leaf_451_CLK _02905_ VGND VGND VPWR VPWR registers\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_237_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_264_CLK clknet_6_60__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_264_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33742_ clknet_leaf_147_CLK _01856_ VGND VGND VPWR VPWR registers\[40\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18676_ registers\[28\]\[8\] registers\[29\]\[8\] registers\[30\]\[8\] registers\[31\]\[8\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__mux4_1
X_30954_ _13965_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__clkbuf_1
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17627_ registers\[48\]\[44\] registers\[49\]\[44\] registers\[50\]\[44\] registers\[51\]\[44\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__mux4_1
XFILLER_58_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33673_ clknet_leaf_245_CLK _01787_ VGND VGND VPWR VPWR registers\[42\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30885_ _13929_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_229_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35412_ clknet_leaf_81_CLK _03526_ VGND VGND VPWR VPWR registers\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32624_ clknet_leaf_367_CLK _00738_ VGND VGND VPWR VPWR registers\[58\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_17558_ _14516_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35343_ clknet_leaf_137_CLK _03457_ VGND VGND VPWR VPWR registers\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16509_ registers\[8\]\[12\] registers\[9\]\[12\] registers\[10\]\[12\] registers\[11\]\[12\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _15011_ sky130_fd_sc_hd__mux4_1
X_32555_ clknet_leaf_401_CLK _00669_ VGND VGND VPWR VPWR registers\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_17489_ _14553_ VGND VGND VPWR VPWR _15963_ sky130_fd_sc_hd__clkbuf_4
XFILLER_220_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_993 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31506_ _09786_ registers\[6\]\[45\] _14250_ VGND VGND VPWR VPWR _14256_ sky130_fd_sc_hd__mux2_1
X_19228_ registers\[8\]\[24\] registers\[9\]\[24\] registers\[10\]\[24\] registers\[11\]\[24\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__mux4_1
X_35274_ clknet_leaf_149_CLK _03388_ VGND VGND VPWR VPWR registers\[17\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32486_ clknet_leaf_451_CLK _00600_ VGND VGND VPWR VPWR registers\[60\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34225_ clknet_leaf_355_CLK _02339_ VGND VGND VPWR VPWR registers\[33\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_31437_ _09683_ registers\[6\]\[12\] _14217_ VGND VGND VPWR VPWR _14220_ sky130_fd_sc_hd__mux2_1
X_19159_ registers\[52\]\[22\] registers\[53\]\[22\] registers\[54\]\[22\] registers\[55\]\[22\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__mux4_1
XFILLER_145_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22170_ _08610_ _08825_ _08826_ _08613_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__a22o_1
X_34156_ clknet_leaf_322_CLK _02270_ VGND VGND VPWR VPWR registers\[34\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31368_ _14183_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33107_ clknet_leaf_70_CLK _01221_ VGND VGND VPWR VPWR registers\[50\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_21121_ registers\[28\]\[12\] registers\[29\]\[12\] registers\[30\]\[12\] registers\[31\]\[12\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__mux4_1
X_30319_ registers\[15\]\[59\] _13058_ _13621_ VGND VGND VPWR VPWR _13631_ sky130_fd_sc_hd__mux2_1
X_34087_ clknet_leaf_431_CLK _02201_ VGND VGND VPWR VPWR registers\[35\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_31299_ _14147_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33038_ clknet_leaf_74_CLK _01152_ VGND VGND VPWR VPWR registers\[51\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21052_ registers\[20\]\[10\] registers\[21\]\[10\] registers\[22\]\[10\] registers\[23\]\[10\]
+ _07739_ _07740_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__mux4_1
XFILLER_232_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _05116_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__buf_4
X_25860_ _10850_ registers\[47\]\[57\] _11214_ VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__mux2_1
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_219_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24811_ _09605_ registers\[54\]\[43\] _10631_ VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__mux2_1
XFILLER_189_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25791_ _10781_ registers\[47\]\[24\] _11181_ VGND VGND VPWR VPWR _11186_ sky130_fd_sc_hd__mux2_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34989_ clknet_leaf_396_CLK _03103_ VGND VGND VPWR VPWR registers\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_255_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_255_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27530_ _11832_ registers\[35\]\[49\] _12122_ VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__mux2_1
X_24742_ _09535_ registers\[54\]\[10\] _10598_ VGND VGND VPWR VPWR _10599_ sky130_fd_sc_hd__mux2_1
XFILLER_55_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ registers\[4\]\[36\] registers\[5\]\[36\] registers\[6\]\[36\] registers\[7\]\[36\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__mux4_1
XFILLER_215_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20905_ registers\[20\]\[6\] registers\[21\]\[6\] registers\[22\]\[6\] registers\[23\]\[6\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__mux4_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27461_ _11763_ registers\[35\]\[16\] _12089_ VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__mux2_1
XFILLER_160_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24673_ _10561_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
X_21885_ registers\[4\]\[34\] registers\[5\]\[34\] registers\[6\]\[34\] registers\[7\]\[34\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__mux4_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29200_ net43 VGND VGND VPWR VPWR _13035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_242_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26412_ _10862_ registers\[43\]\[63\] _11442_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__mux2_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _07386_ _07529_ _07530_ _07396_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__a22o_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _09974_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27392_ _12059_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29131_ _12988_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26343_ _11442_ VGND VGND VPWR VPWR _11476_ sky130_fd_sc_hd__clkbuf_8
X_23555_ _09642_ registers\[19\]\[61\] _09869_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__mux2_1
X_20767_ _07388_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__buf_6
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22506_ _07285_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__buf_4
XFILLER_211_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_210_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29062_ registers\[23\]\[3\] _12941_ _12935_ VGND VGND VPWR VPWR _12942_ sky130_fd_sc_hd__mux2_1
X_26274_ _11439_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
X_23486_ _09573_ registers\[19\]\[28\] _09892_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__mux2_1
X_20698_ _07386_ _07390_ _07394_ _07396_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__a22o_1
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28013_ _12387_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22437_ registers\[48\]\[50\] registers\[49\]\[50\] registers\[50\]\[50\] registers\[51\]\[50\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__mux4_1
XFILLER_108_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25225_ _10883_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25156_ net49 VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__clkbuf_4
X_22368_ _09012_ _09014_ _09017_ _09018_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__a22o_1
XFILLER_191_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_237_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24107_ _10230_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
X_21319_ _07924_ _07998_ _07999_ _07927_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__a22o_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25087_ _10795_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
X_29964_ _13444_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__clkbuf_1
X_22299_ _08946_ _08951_ _08748_ _08749_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__o211a_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28915_ registers\[24\]\[0\] _10303_ _12861_ VGND VGND VPWR VPWR _12862_ sky130_fd_sc_hd__mux2_1
X_24038_ _09577_ registers\[5\]\[30\] _10194_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__mux2_1
X_29895_ _13352_ VGND VGND VPWR VPWR _13408_ sky130_fd_sc_hd__buf_4
XFILLER_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_984 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28846_ _12825_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__clkbuf_1
X_16860_ _15206_ _15350_ _15351_ _15210_ VGND VGND VPWR VPWR _15352_ sky130_fd_sc_hd__a22o_1
XFILLER_215_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_219_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28777_ _12788_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__clkbuf_1
X_16791_ registers\[12\]\[20\] registers\[13\]\[20\] registers\[14\]\[20\] registers\[15\]\[20\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15285_ sky130_fd_sc_hd__mux4_1
XFILLER_92_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25989_ _10844_ registers\[46\]\[54\] _11285_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_246_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_246_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_234_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18530_ _05113_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__buf_4
XFILLER_19_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27728_ _12237_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__clkbuf_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _05119_ _05220_ _05221_ _05131_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__a22o_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27659_ registers\[34\]\[45\] _10399_ _12195_ VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__mux2_1
XFILLER_45_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_241 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_252 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _14543_ VGND VGND VPWR VPWR _15888_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_263 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18392_ _05079_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__buf_4
XFILLER_18_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30670_ _13816_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__clkbuf_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_296 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29329_ _13110_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_38__f_CLK clknet_5_19_0_CLK VGND VGND VPWR VPWR clknet_6_38__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_17343_ _14548_ VGND VGND VPWR VPWR _15821_ sky130_fd_sc_hd__buf_4
XFILLER_14_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32340_ clknet_leaf_64_CLK _00454_ VGND VGND VPWR VPWR registers\[61\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17274_ registers\[48\]\[34\] registers\[49\]\[34\] registers\[50\]\[34\] registers\[51\]\[34\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15754_ sky130_fd_sc_hd__mux4_1
XFILLER_9_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19013_ registers\[52\]\[18\] registers\[53\]\[18\] registers\[54\]\[18\] registers\[55\]\[18\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__mux4_1
X_16225_ registers\[12\]\[4\] registers\[13\]\[4\] registers\[14\]\[4\] registers\[15\]\[4\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14735_ sky130_fd_sc_hd__mux4_1
XFILLER_158_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32271_ clknet_leaf_113_CLK _00385_ VGND VGND VPWR VPWR registers\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34010_ clknet_leaf_25_CLK _02124_ VGND VGND VPWR VPWR registers\[36\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_31222_ _14106_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__clkbuf_1
X_16156_ registers\[8\]\[2\] registers\[9\]\[2\] registers\[10\]\[2\] registers\[11\]\[2\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _14668_ sky130_fd_sc_hd__mux4_1
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31153_ _14070_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__clkbuf_1
X_16087_ _14600_ VGND VGND VPWR VPWR _14601_ sky130_fd_sc_hd__buf_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30104_ _13518_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__clkbuf_1
X_19915_ _06631_ _06634_ _06537_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__o21ba_1
XFILLER_29_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35961_ clknet_leaf_315_CLK _04075_ VGND VGND VPWR VPWR registers\[6\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_31084_ registers\[0\]\[37\] _13012_ _14026_ VGND VGND VPWR VPWR _14034_ sky130_fd_sc_hd__mux2_1
XFILLER_69_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_485_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_485_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_30035_ registers\[17\]\[52\] _13044_ _13479_ VGND VGND VPWR VPWR _13482_ sky130_fd_sc_hd__mux2_1
X_34912_ clknet_leaf_490_CLK _03026_ VGND VGND VPWR VPWR registers\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19846_ _06546_ _06553_ _06560_ _06567_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__or4_4
XFILLER_110_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35892_ clknet_leaf_418_CLK _04006_ VGND VGND VPWR VPWR registers\[7\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_110_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34843_ clknet_leaf_490_CLK _02957_ VGND VGND VPWR VPWR registers\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19777_ _05097_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__clkbuf_4
X_16989_ _14546_ VGND VGND VPWR VPWR _15477_ sky130_fd_sc_hd__buf_6
XFILLER_84_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_237_CLK clknet_6_61__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_237_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18728_ registers\[52\]\[10\] registers\[53\]\[10\] registers\[54\]\[10\] registers\[55\]\[10\]
+ _05340_ _05341_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux4_1
X_34774_ clknet_leaf_87_CLK _02888_ VGND VGND VPWR VPWR registers\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_31986_ clknet_leaf_22_CLK _00157_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_225_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33725_ clknet_leaf_278_CLK _01839_ VGND VGND VPWR VPWR registers\[41\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_18659_ registers\[60\]\[8\] registers\[61\]\[8\] registers\[62\]\[8\] registers\[63\]\[8\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__mux4_1
X_30937_ registers\[10\]\[31\] _13000_ _13955_ VGND VGND VPWR VPWR _13957_ sky130_fd_sc_hd__mux2_1
XFILLER_224_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21670_ registers\[8\]\[28\] registers\[9\]\[28\] registers\[10\]\[28\] registers\[11\]\[28\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__mux4_1
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30868_ _09825_ registers\[11\]\[63\] _13850_ VGND VGND VPWR VPWR _13920_ sky130_fd_sc_hd__mux2_1
X_33656_ clknet_leaf_338_CLK _01770_ VGND VGND VPWR VPWR registers\[42\]\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20621_ _07281_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32607_ clknet_leaf_38_CLK _00721_ VGND VGND VPWR VPWR registers\[58\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33587_ clknet_leaf_348_CLK _01701_ VGND VGND VPWR VPWR registers\[43\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30799_ _13850_ VGND VGND VPWR VPWR _13884_ sky130_fd_sc_hd__buf_4
XFILLER_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23340_ registers\[9\]\[61\] _09821_ _09708_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__mux2_1
XFILLER_123_1316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20552_ registers\[56\]\[63\] registers\[57\]\[63\] registers\[58\]\[63\] registers\[59\]\[63\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__mux4_1
X_35326_ clknet_leaf_191_CLK _03440_ VGND VGND VPWR VPWR registers\[16\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_32538_ clknet_leaf_475_CLK _00652_ VGND VGND VPWR VPWR registers\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23271_ _09708_ VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__buf_4
X_20483_ _07164_ _07171_ _07178_ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__or4_1
X_32469_ clknet_leaf_182_CLK _00583_ VGND VGND VPWR VPWR registers\[60\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_35257_ clknet_leaf_309_CLK _03371_ VGND VGND VPWR VPWR registers\[17\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25010_ net61 VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__buf_4
X_22222_ registers\[36\]\[44\] registers\[37\]\[44\] registers\[38\]\[44\] registers\[39\]\[44\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__mux4_1
X_34208_ clknet_leaf_17_CLK _02322_ VGND VGND VPWR VPWR registers\[33\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35188_ clknet_leaf_417_CLK _03302_ VGND VGND VPWR VPWR registers\[18\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22153_ _07285_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__clkbuf_4
X_34139_ clknet_leaf_18_CLK _02253_ VGND VGND VPWR VPWR registers\[34\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21104_ _07640_ _07789_ _07790_ _07646_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__a22o_1
XTAP_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26961_ _11823_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22084_ registers\[48\]\[40\] registers\[49\]\[40\] registers\[50\]\[40\] registers\[51\]\[40\]
+ _08672_ _08673_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__mux4_1
XTAP_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_476_CLK clknet_6_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_476_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28700_ _12748_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25912_ _11249_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
X_21035_ _07349_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29680_ _13295_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__clkbuf_1
X_26892_ _11776_ registers\[3\]\[22\] _11772_ VGND VGND VPWR VPWR _11777_ sky130_fd_sc_hd__mux2_1
XFILLER_248_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28631_ _11851_ registers\[27\]\[58\] _12703_ VGND VGND VPWR VPWR _12712_ sky130_fd_sc_hd__mux2_1
XFILLER_219_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25843_ _10833_ registers\[47\]\[49\] _11203_ VGND VGND VPWR VPWR _11213_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_228_CLK clknet_6_55__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_228_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28562_ _11782_ registers\[27\]\[25\] _12670_ VGND VGND VPWR VPWR _12676_ sky130_fd_sc_hd__mux2_1
X_25774_ _10764_ registers\[47\]\[16\] _11170_ VGND VGND VPWR VPWR _11177_ sky130_fd_sc_hd__mux2_1
X_22986_ _09586_ registers\[62\]\[34\] _09578_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__mux2_1
XFILLER_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27513_ _12123_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24725_ _09519_ registers\[54\]\[2\] _10587_ VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__mux2_1
XFILLER_243_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28493_ _12639_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__clkbuf_1
X_21937_ _08596_ _08599_ _08397_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__o21ba_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27444_ _11746_ registers\[35\]\[8\] _12078_ VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__mux2_1
XFILLER_203_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24656_ _10552_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21868_ registers\[44\]\[34\] registers\[45\]\[34\] registers\[46\]\[34\] registers\[47\]\[34\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__mux4_1
XFILLER_169_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ registers\[61\]\[20\] _09699_ _09965_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__mux2_1
X_20819_ registers\[52\]\[4\] registers\[53\]\[4\] registers\[54\]\[4\] registers\[55\]\[4\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__mux4_1
X_27375_ _12050_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24587_ _10516_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21799_ registers\[32\]\[32\] registers\[33\]\[32\] registers\[34\]\[32\] registers\[35\]\[32\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__mux4_1
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_400_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_400_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_29114_ _12934_ VGND VGND VPWR VPWR _12977_ sky130_fd_sc_hd__buf_4
XFILLER_184_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26326_ _11467_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_1
X_23538_ _09928_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29045_ _12929_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__clkbuf_1
X_26257_ _10842_ registers\[44\]\[53\] _11427_ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__mux2_1
XFILLER_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23469_ _09869_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__buf_4
X_16010_ net69 net70 VGND VGND VPWR VPWR _14524_ sky130_fd_sc_hd__or2b_4
XFILLER_137_862 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25208_ _10874_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26188_ _10772_ registers\[44\]\[20\] _11394_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__mux2_1
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25139_ _10830_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _04729_ _04734_ _04630_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__o21ba_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29947_ registers\[17\]\[10\] _12955_ _13435_ VGND VGND VPWR VPWR _13436_ sky130_fd_sc_hd__mux2_1
XFILLER_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19700_ _06425_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_467_CLK clknet_6_8__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_467_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16912_ registers\[40\]\[24\] registers\[41\]\[24\] registers\[42\]\[24\] registers\[43\]\[24\]
+ _15335_ _15336_ VGND VGND VPWR VPWR _15402_ sky130_fd_sc_hd__mux4_1
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17892_ registers\[24\]\[51\] registers\[25\]\[51\] registers\[26\]\[51\] registers\[27\]\[51\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__mux4_1
X_29878_ _13399_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19631_ registers\[40\]\[36\] registers\[41\]\[36\] registers\[42\]\[36\] registers\[43\]\[36\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__mux4_1
X_16843_ _14493_ VGND VGND VPWR VPWR _15335_ sky130_fd_sc_hd__buf_4
X_28829_ _12816_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_219_CLK clknet_6_53__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_219_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31840_ _09681_ registers\[49\]\[11\] _14430_ VGND VGND VPWR VPWR _14432_ sky130_fd_sc_hd__mux2_1
X_19562_ _06288_ _06291_ _06194_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__o21ba_1
XFILLER_93_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16774_ _14998_ _15266_ _15267_ _15001_ VGND VGND VPWR VPWR _15268_ sky130_fd_sc_hd__a22o_1
XFILLER_225_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_234_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18513_ _05078_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__buf_6
XFILLER_218_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31771_ _14395_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__clkbuf_1
X_19493_ _06203_ _06210_ _06217_ _06224_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__or4_1
XFILLER_222_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ registers\[44\]\[2\] registers\[45\]\[2\] registers\[46\]\[2\] registers\[47\]\[2\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__mux4_1
X_30722_ _13843_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__clkbuf_1
X_33510_ clknet_leaf_60_CLK _01624_ VGND VGND VPWR VPWR registers\[44\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34490_ clknet_leaf_302_CLK _02604_ VGND VGND VPWR VPWR registers\[2\]\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33441_ clknet_leaf_35_CLK _01555_ VGND VGND VPWR VPWR registers\[45\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_18375_ _05125_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__buf_6
X_30653_ _13807_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__clkbuf_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1081 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17326_ registers\[20\]\[35\] registers\[21\]\[35\] registers\[22\]\[35\] registers\[23\]\[35\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15805_ sky130_fd_sc_hd__mux4_1
X_36160_ clknet_leaf_270_CLK _04274_ VGND VGND VPWR VPWR registers\[49\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_33372_ clknet_leaf_29_CLK _01486_ VGND VGND VPWR VPWR registers\[46\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_30584_ _09810_ registers\[13\]\[56\] _13764_ VGND VGND VPWR VPWR _13771_ sky130_fd_sc_hd__mux2_1
XFILLER_175_935 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32323_ clknet_leaf_221_CLK _00437_ VGND VGND VPWR VPWR registers\[19\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_35111_ clknet_leaf_463_CLK _03225_ VGND VGND VPWR VPWR registers\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_36091_ clknet_leaf_284_CLK _04205_ VGND VGND VPWR VPWR registers\[59\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_17257_ registers\[16\]\[33\] registers\[17\]\[33\] registers\[18\]\[33\] registers\[19\]\[33\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15738_ sky130_fd_sc_hd__mux4_1
XFILLER_70_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16208_ _14648_ _14716_ _14717_ _14653_ VGND VGND VPWR VPWR _14718_ sky130_fd_sc_hd__a22o_1
X_35042_ clknet_leaf_471_CLK _03156_ VGND VGND VPWR VPWR registers\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_32254_ clknet_leaf_268_CLK _00368_ VGND VGND VPWR VPWR registers\[39\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17188_ _15633_ _15669_ _15670_ _15636_ VGND VGND VPWR VPWR _15671_ sky130_fd_sc_hd__a22o_1
XFILLER_157_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31205_ registers\[8\]\[30\] net24 _14097_ VGND VGND VPWR VPWR _14098_ sky130_fd_sc_hd__mux2_1
X_16139_ registers\[40\]\[2\] registers\[41\]\[2\] registers\[42\]\[2\] registers\[43\]\[2\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14651_ sky130_fd_sc_hd__mux4_1
XFILLER_192_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32185_ clknet_leaf_484_CLK _00299_ VGND VGND VPWR VPWR registers\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31136_ registers\[0\]\[62\] _13064_ _13992_ VGND VGND VPWR VPWR _14061_ sky130_fd_sc_hd__mux2_1
XFILLER_143_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_458_CLK clknet_6_10__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_458_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35944_ clknet_leaf_400_CLK _04058_ VGND VGND VPWR VPWR registers\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_31067_ registers\[0\]\[29\] _12995_ _14015_ VGND VGND VPWR VPWR _14025_ sky130_fd_sc_hd__mux2_1
X_30018_ registers\[17\]\[44\] _13027_ _13468_ VGND VGND VPWR VPWR _13473_ sky130_fd_sc_hd__mux2_1
XFILLER_5_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19829_ registers\[52\]\[41\] registers\[53\]\[41\] registers\[54\]\[41\] registers\[55\]\[41\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__mux4_1
XFILLER_233_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35875_ clknet_leaf_470_CLK _03989_ VGND VGND VPWR VPWR registers\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34826_ clknet_leaf_153_CLK _02940_ VGND VGND VPWR VPWR registers\[24\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22840_ registers\[20\]\[62\] registers\[21\]\[62\] registers\[22\]\[62\] registers\[23\]\[62\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__mux4_1
XFILLER_83_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34757_ clknet_leaf_219_CLK _02871_ VGND VGND VPWR VPWR registers\[25\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_22771_ _07276_ _09408_ _09409_ _07286_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__a22o_1
XFILLER_25_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31969_ clknet_leaf_5_CLK _00138_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24510_ _10474_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_227_1137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21722_ _08119_ _08389_ _08390_ _08124_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__a22o_1
X_33708_ clknet_leaf_326_CLK _01822_ VGND VGND VPWR VPWR registers\[41\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_25490_ _11025_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34688_ clknet_leaf_222_CLK _02802_ VGND VGND VPWR VPWR registers\[26\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24441_ registers\[57\]\[63\] _10436_ net283 VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__mux2_1
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21653_ _08126_ _08322_ _08323_ _08129_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__a22o_1
X_33639_ clknet_leaf_430_CLK _01753_ VGND VGND VPWR VPWR registers\[42\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_21__f_CLK clknet_5_10_0_CLK VGND VGND VPWR VPWR clknet_6_21__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_27160_ _11732_ registers\[37\]\[1\] _11936_ VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__mux2_1
X_20604_ _07277_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__buf_12
XFILLER_162_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21584_ _08253_ _08256_ _08054_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__o21ba_1
X_24372_ _10390_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26111_ _10831_ registers\[45\]\[48\] _11345_ VGND VGND VPWR VPWR _11354_ sky130_fd_sc_hd__mux2_1
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23323_ registers\[9\]\[56\] _09810_ _09798_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__mux2_1
X_20535_ _07232_ _07235_ _05133_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__o21ba_1
X_35309_ clknet_leaf_397_CLK _03423_ VGND VGND VPWR VPWR registers\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_27091_ _11901_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26042_ _10762_ registers\[45\]\[15\] _11312_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__mux2_1
X_20466_ registers\[52\]\[60\] registers\[53\]\[60\] registers\[54\]\[60\] registers\[55\]\[60\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__mux4_1
XFILLER_14_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23254_ registers\[9\]\[35\] _09764_ _09754_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__mux2_1
XFILLER_165_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22205_ registers\[12\]\[43\] registers\[13\]\[43\] registers\[14\]\[43\] registers\[15\]\[43\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__mux4_1
XFILLER_101_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23185_ registers\[9\]\[10\] _09678_ _09722_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__mux2_1
XFILLER_238_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20397_ _06912_ _07100_ _07101_ _06917_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__a22o_1
XTAP_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29801_ registers\[18\]\[5\] _12945_ _13353_ VGND VGND VPWR VPWR _13359_ sky130_fd_sc_hd__mux2_1
X_22136_ registers\[4\]\[41\] registers\[5\]\[41\] registers\[6\]\[41\] registers\[7\]\[41\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__mux4_1
XTAP_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1409 _00179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27993_ _11753_ registers\[31\]\[11\] _12375_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__mux2_1
Xoutput270 net270 VGND VGND VPWR VPWR D3[57] sky130_fd_sc_hd__buf_2
XTAP_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput281 net281 VGND VGND VPWR VPWR D3[9] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_449_CLK clknet_6_11__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_449_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29732_ _13322_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__clkbuf_1
X_22067_ registers\[28\]\[39\] registers\[29\]\[39\] registers\[30\]\[39\] registers\[31\]\[39\]
+ _08492_ _08493_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__mux4_1
X_26944_ _11811_ registers\[3\]\[39\] _11793_ VGND VGND VPWR VPWR _11812_ sky130_fd_sc_hd__mux2_1
XFILLER_248_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21018_ _07289_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29663_ _13286_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26875_ net9 VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__clkbuf_4
XTAP_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28614_ _12647_ VGND VGND VPWR VPWR _12703_ sky130_fd_sc_hd__buf_4
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25826_ _11204_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
X_29594_ registers\[20\]\[35\] _13008_ _13244_ VGND VGND VPWR VPWR _13250_ sky130_fd_sc_hd__mux2_1
XFILLER_235_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28545_ _11765_ registers\[27\]\[17\] _12659_ VGND VGND VPWR VPWR _12667_ sky130_fd_sc_hd__mux2_1
X_25757_ _10747_ registers\[47\]\[8\] _11159_ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__mux2_1
XFILLER_204_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22969_ net22 VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__buf_2
XFILLER_245_1204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24708_ _10579_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28476_ _12630_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__clkbuf_1
X_16490_ _14493_ VGND VGND VPWR VPWR _14992_ sky130_fd_sc_hd__buf_4
XFILLER_167_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25688_ registers\[48\]\[40\] _10388_ _11130_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__mux2_1
XFILLER_215_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27427_ _12077_ VGND VGND VPWR VPWR _12078_ sky130_fd_sc_hd__buf_6
X_24639_ _10543_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18160_ _04683_ _04925_ _04926_ _04686_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__a22o_1
XFILLER_141_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27358_ registers\[36\]\[31\] _10370_ _12040_ VGND VGND VPWR VPWR _12042_ sky130_fd_sc_hd__mux2_1
X_17111_ registers\[24\]\[29\] registers\[25\]\[29\] registers\[26\]\[29\] registers\[27\]\[29\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15596_ sky130_fd_sc_hd__mux4_1
XFILLER_129_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26309_ _11458_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
X_18091_ _04637_ _04859_ _04860_ _04642_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__a22o_1
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27289_ _11861_ registers\[37\]\[63\] _11935_ VGND VGND VPWR VPWR _12005_ sky130_fd_sc_hd__mux2_1
XFILLER_172_905 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29028_ registers\[24\]\[54\] _10418_ _12916_ VGND VGND VPWR VPWR _12921_ sky130_fd_sc_hd__mux2_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17042_ registers\[28\]\[27\] registers\[29\]\[27\] registers\[30\]\[27\] registers\[31\]\[27\]
+ _15364_ _15365_ VGND VGND VPWR VPWR _15529_ sky130_fd_sc_hd__mux4_1
XFILLER_125_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18993_ _05717_ _05724_ _05731_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__or4_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17944_ _04683_ _04716_ _04717_ _04686_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a22o_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33990_ clknet_leaf_246_CLK _02104_ VGND VGND VPWR VPWR registers\[37\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17875_ registers\[36\]\[51\] registers\[37\]\[51\] registers\[38\]\[51\] registers\[39\]\[51\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__mux4_1
X_32941_ clknet_leaf_373_CLK _01055_ VGND VGND VPWR VPWR registers\[53\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19614_ _05053_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__buf_4
X_35660_ clknet_leaf_144_CLK _03774_ VGND VGND VPWR VPWR registers\[11\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_16826_ registers\[8\]\[21\] registers\[9\]\[21\] registers\[10\]\[21\] registers\[11\]\[21\]
+ _15106_ _15107_ VGND VGND VPWR VPWR _15319_ sky130_fd_sc_hd__mux4_1
XFILLER_94_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32872_ clknet_leaf_423_CLK _00986_ VGND VGND VPWR VPWR registers\[54\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34611_ clknet_leaf_408_CLK _02725_ VGND VGND VPWR VPWR registers\[27\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_31823_ _09664_ registers\[49\]\[3\] _14419_ VGND VGND VPWR VPWR _14423_ sky130_fd_sc_hd__mux2_1
X_16757_ _15248_ _15251_ _14945_ VGND VGND VPWR VPWR _15252_ sky130_fd_sc_hd__o21ba_1
X_19545_ _06098_ _06273_ _06274_ _06102_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__a22o_1
X_35591_ clknet_leaf_214_CLK _03705_ VGND VGND VPWR VPWR registers\[12\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31754_ _14386_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__clkbuf_1
X_34542_ clknet_leaf_387_CLK _02656_ VGND VGND VPWR VPWR registers\[28\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_19476_ registers\[52\]\[31\] registers\[53\]\[31\] registers\[54\]\[31\] registers\[55\]\[31\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__mux4_1
X_16688_ _14947_ _15183_ _15184_ _14950_ VGND VGND VPWR VPWR _15185_ sky130_fd_sc_hd__a22o_1
XFILLER_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30705_ _13834_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_222_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18427_ registers\[24\]\[1\] registers\[25\]\[1\] registers\[26\]\[1\] registers\[27\]\[1\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__mux4_1
XFILLER_72_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31685_ _14350_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__clkbuf_1
X_34473_ clknet_leaf_458_CLK _02587_ VGND VGND VPWR VPWR registers\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36212_ clknet_leaf_115_CLK _00095_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dfxtp_1
XFILLER_166_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33424_ clknet_leaf_129_CLK _01538_ VGND VGND VPWR VPWR registers\[45\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_18358_ _05120_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__buf_8
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30636_ _13798_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_5_19_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_19_0_CLK sky130_fd_sc_hd__clkbuf_8
X_17309_ registers\[60\]\[35\] registers\[61\]\[35\] registers\[62\]\[35\] registers\[63\]\[35\]
+ _15756_ _15550_ VGND VGND VPWR VPWR _15788_ sky130_fd_sc_hd__mux4_1
X_33355_ clknet_leaf_165_CLK _01469_ VGND VGND VPWR VPWR registers\[47\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_36143_ clknet_leaf_365_CLK _04257_ VGND VGND VPWR VPWR registers\[49\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_18289_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__buf_4
XFILLER_175_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30567_ _09793_ registers\[13\]\[48\] _13753_ VGND VGND VPWR VPWR _13762_ sky130_fd_sc_hd__mux2_1
XFILLER_30_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20320_ registers\[0\]\[55\] registers\[1\]\[55\] registers\[2\]\[55\] registers\[3\]\[55\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__mux4_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32306_ clknet_leaf_412_CLK _00420_ VGND VGND VPWR VPWR registers\[19\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_33286_ clknet_leaf_261_CLK _01400_ VGND VGND VPWR VPWR registers\[48\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_36074_ clknet_leaf_420_CLK _04188_ VGND VGND VPWR VPWR registers\[59\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_30498_ _09689_ registers\[13\]\[15\] _13720_ VGND VGND VPWR VPWR _13726_ sky130_fd_sc_hd__mux2_1
X_35025_ clknet_leaf_113_CLK _03139_ VGND VGND VPWR VPWR registers\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_20251_ _06784_ _06959_ _06960_ _06788_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__a22o_1
X_32237_ clknet_leaf_327_CLK _00351_ VGND VGND VPWR VPWR registers\[39\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_1111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20182_ registers\[52\]\[51\] registers\[53\]\[51\] registers\[54\]\[51\] registers\[55\]\[51\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__mux4_1
X_32168_ clknet_leaf_106_CLK _00282_ VGND VGND VPWR VPWR registers\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31119_ _14052_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24990_ _09941_ _10584_ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__nor2_8
X_32099_ clknet_leaf_483_CLK _00013_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dfxtp_1
XFILLER_215_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23941_ _09617_ registers\[60\]\[49\] _10133_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__mux2_1
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35927_ clknet_leaf_83_CLK _04041_ VGND VGND VPWR VPWR registers\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26660_ _11643_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__clkbuf_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35858_ clknet_leaf_76_CLK _03972_ VGND VGND VPWR VPWR registers\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23872_ _09548_ registers\[60\]\[16\] _10100_ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__mux2_1
XFILLER_151_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25611_ _11090_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
X_22823_ registers\[48\]\[62\] registers\[49\]\[62\] registers\[50\]\[62\] registers\[51\]\[62\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__mux4_1
XANTENNA_807 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34809_ clknet_leaf_314_CLK _02923_ VGND VGND VPWR VPWR registers\[24\]\[43\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_818 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26591_ _10770_ registers\[41\]\[19\] _11597_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__mux2_1
X_35789_ clknet_leaf_148_CLK _03903_ VGND VGND VPWR VPWR registers\[0\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_232_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_829 _09147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28330_ registers\[2\]\[43\] _10395_ _12550_ VGND VGND VPWR VPWR _12554_ sky130_fd_sc_hd__mux2_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25542_ _11052_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__clkbuf_1
X_22754_ _09393_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21705_ registers\[0\]\[29\] registers\[1\]\[29\] registers\[2\]\[29\] registers\[3\]\[29\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__mux4_1
X_28261_ registers\[2\]\[10\] _10325_ _12517_ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__mux2_1
X_25473_ _11016_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_1
X_22685_ _09323_ _09326_ _09102_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__o21ba_1
XFILLER_212_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27212_ _11784_ registers\[37\]\[26\] _11958_ VGND VGND VPWR VPWR _11965_ sky130_fd_sc_hd__mux2_1
X_24424_ _10425_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
X_21636_ registers\[4\]\[27\] registers\[5\]\[27\] registers\[6\]\[27\] registers\[7\]\[27\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__mux4_1
X_28192_ _12481_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27143_ _11928_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24355_ registers\[57\]\[35\] _10378_ _10368_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__mux2_1
X_21567_ _07929_ _08239_ _08240_ _07932_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__a22o_1
XFILLER_60_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23306_ _09799_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20518_ registers\[44\]\[62\] registers\[45\]\[62\] registers\[46\]\[62\] registers\[47\]\[62\]
+ _05096_ _05098_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__mux4_1
XFILLER_125_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27074_ _11892_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21498_ _07305_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__buf_4
X_24286_ net5 VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__buf_4
XFILLER_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26025_ _10745_ registers\[45\]\[7\] _11301_ VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__mux2_1
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20449_ registers\[28\]\[59\] registers\[29\]\[59\] registers\[30\]\[59\] registers\[31\]\[59\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__mux4_1
XFILLER_181_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23237_ net24 VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_865 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23168_ _09713_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
XTAP_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1206 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1217 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1228 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22119_ registers\[32\]\[41\] registers\[33\]\[41\] registers\[34\]\[41\] registers\[35\]\[41\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__mux4_1
X_15990_ _14495_ VGND VGND VPWR VPWR _14504_ sky130_fd_sc_hd__buf_12
XTAP_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27976_ _11736_ registers\[31\]\[3\] _12364_ VGND VGND VPWR VPWR _12368_ sky130_fd_sc_hd__mux2_1
X_23099_ net45 VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__buf_4
XANTENNA_1239 _00088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26927_ _11800_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_1
X_29715_ _13313_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__clkbuf_1
XTAP_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ registers\[48\]\[45\] registers\[49\]\[45\] registers\[50\]\[45\] registers\[51\]\[45\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__mux4_1
X_29646_ registers\[20\]\[60\] _13060_ _13210_ VGND VGND VPWR VPWR _13277_ sky130_fd_sc_hd__mux2_1
XTAP_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26858_ _11753_ registers\[3\]\[11\] _11751_ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__mux2_1
XFILLER_76_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16611_ _14796_ _15108_ _15109_ _14799_ VGND VGND VPWR VPWR _15110_ sky130_fd_sc_hd__a22o_1
XFILLER_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_882 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25809_ _11195_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17591_ _04340_ _04373_ _04374_ _04343_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a22o_1
XFILLER_112_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29577_ registers\[20\]\[27\] _12991_ _13233_ VGND VGND VPWR VPWR _13241_ sky130_fd_sc_hd__mux2_1
XFILLER_91_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26789_ _11711_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28528_ _11748_ registers\[27\]\[9\] _12648_ VGND VGND VPWR VPWR _12658_ sky130_fd_sc_hd__mux2_1
X_16542_ registers\[0\]\[13\] registers\[1\]\[13\] registers\[2\]\[13\] registers\[3\]\[13\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15043_ sky130_fd_sc_hd__mux4_1
X_19330_ _05755_ _06064_ _06065_ _05759_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__a22o_1
XFILLER_56_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19261_ _05053_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__buf_4
XFILLER_95_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16473_ registers\[8\]\[11\] registers\[9\]\[11\] registers\[10\]\[11\] registers\[11\]\[11\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _14976_ sky130_fd_sc_hd__mux4_1
X_28459_ _11813_ registers\[28\]\[40\] _12621_ VGND VGND VPWR VPWR _12622_ sky130_fd_sc_hd__mux2_1
X_18212_ _04974_ _04977_ _14613_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__o21ba_1
X_31470_ _09749_ registers\[6\]\[28\] _14228_ VGND VGND VPWR VPWR _14237_ sky130_fd_sc_hd__mux2_1
X_19192_ _05755_ _05930_ _05931_ _05759_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__a22o_1
XFILLER_223_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18143_ registers\[4\]\[59\] registers\[5\]\[59\] registers\[6\]\[59\] registers\[7\]\[59\]
+ _14589_ _14590_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__mux4_1
X_30421_ _13685_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33140_ clknet_leaf_350_CLK _01254_ VGND VGND VPWR VPWR registers\[50\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_18074_ _04540_ _04842_ _04843_ _04546_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a22o_1
X_30352_ _13637_ VGND VGND VPWR VPWR _13649_ sky130_fd_sc_hd__buf_4
XFILLER_171_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17025_ registers\[56\]\[27\] registers\[57\]\[27\] registers\[58\]\[27\] registers\[59\]\[27\]
+ _15409_ _15199_ VGND VGND VPWR VPWR _15512_ sky130_fd_sc_hd__mux4_1
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33071_ clknet_leaf_364_CLK _01185_ VGND VGND VPWR VPWR registers\[51\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30283_ _13612_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__clkbuf_1
X_32022_ clknet_leaf_66_CLK _00200_ VGND VGND VPWR VPWR registers\[62\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ registers\[52\]\[17\] registers\[53\]\[17\] registers\[54\]\[17\] registers\[55\]\[17\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__mux4_1
XFILLER_234_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1740 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1751 _06911_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _04698_ _04701_ _04630_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__o21ba_1
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_1225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1762 _07392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1773 _11371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33973_ clknet_leaf_350_CLK _02087_ VGND VGND VPWR VPWR registers\[37\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1784 _14518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35712_ clknet_leaf_240_CLK _03826_ VGND VGND VPWR VPWR registers\[10\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_32924_ clknet_leaf_53_CLK _01038_ VGND VGND VPWR VPWR registers\[53\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_17858_ _14567_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35643_ clknet_leaf_300_CLK _03757_ VGND VGND VPWR VPWR registers\[11\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_16809_ _15294_ _15301_ _15302_ VGND VGND VPWR VPWR _15303_ sky130_fd_sc_hd__o21ba_1
X_32855_ clknet_leaf_62_CLK _00969_ VGND VGND VPWR VPWR registers\[54\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_214_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17789_ registers\[20\]\[48\] registers\[21\]\[48\] registers\[22\]\[48\] registers\[23\]\[48\]
+ _04296_ _04297_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__mux4_1
XFILLER_223_931 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31806_ _14413_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__clkbuf_1
X_19528_ registers\[20\]\[32\] registers\[21\]\[32\] registers\[22\]\[32\] registers\[23\]\[32\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux4_1
XFILLER_35_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35574_ clknet_leaf_321_CLK _03688_ VGND VGND VPWR VPWR registers\[12\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_32786_ clknet_leaf_174_CLK _00900_ VGND VGND VPWR VPWR registers\[55\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_2_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_2_0_CLK sky130_fd_sc_hd__clkbuf_8
X_34525_ clknet_leaf_492_CLK _02639_ VGND VGND VPWR VPWR registers\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19459_ _05159_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__clkbuf_4
X_31737_ _14377_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22470_ _09118_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
X_34456_ clknet_leaf_11_CLK _02570_ VGND VGND VPWR VPWR registers\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_31668_ registers\[63\]\[58\] net54 _14332_ VGND VGND VPWR VPWR _14341_ sky130_fd_sc_hd__mux2_1
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33407_ clknet_leaf_273_CLK _01521_ VGND VGND VPWR VPWR registers\[46\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21421_ _07983_ _08097_ _08098_ _07989_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__a22o_1
XFILLER_202_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30619_ _13789_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34387_ clknet_leaf_102_CLK _02501_ VGND VGND VPWR VPWR registers\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31599_ registers\[63\]\[25\] net18 _14299_ VGND VGND VPWR VPWR _14305_ sky130_fd_sc_hd__mux2_1
XFILLER_120_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21352_ registers\[0\]\[19\] registers\[1\]\[19\] registers\[2\]\[19\] registers\[3\]\[19\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__mux4_1
X_24140_ _09544_ registers\[58\]\[14\] _10244_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__mux2_1
X_36126_ clknet_leaf_37_CLK _04240_ VGND VGND VPWR VPWR registers\[49\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_33338_ clknet_leaf_279_CLK _01452_ VGND VGND VPWR VPWR registers\[47\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20303_ _06986_ _06995_ _07002_ _07011_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__or4_4
XFILLER_198_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24071_ _09611_ registers\[5\]\[46\] _10205_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__mux2_1
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36057_ clknet_leaf_84_CLK _04171_ VGND VGND VPWR VPWR registers\[59\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_21283_ registers\[4\]\[17\] registers\[5\]\[17\] registers\[6\]\[17\] registers\[7\]\[17\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__mux4_1
XFILLER_146_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33269_ clknet_leaf_350_CLK _01383_ VGND VGND VPWR VPWR registers\[48\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_20234_ registers\[20\]\[52\] registers\[21\]\[52\] registers\[22\]\[52\] registers\[23\]\[52\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__mux4_1
X_35008_ clknet_leaf_203_CLK _03122_ VGND VGND VPWR VPWR registers\[21\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_23022_ net41 VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1050 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27830_ _12290_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20165_ _05130_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__clkbuf_4
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27761_ _12254_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__clkbuf_1
X_20096_ _05053_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__buf_4
X_24973_ _09632_ registers\[53\]\[56\] _10713_ VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__mux2_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_944 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29500_ _13200_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__clkbuf_1
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26712_ _11671_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23924_ _10134_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
X_27692_ registers\[34\]\[61\] _10432_ _12150_ VGND VGND VPWR VPWR _12218_ sky130_fd_sc_hd__mux2_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29431_ _13164_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26643_ _11634_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _09531_ registers\[60\]\[8\] _10089_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__mux2_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_604 _05097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_615 _05113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_626 _05121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_22806_ registers\[24\]\[61\] registers\[25\]\[61\] registers\[26\]\[61\] registers\[27\]\[61\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__mux4_1
X_29362_ _09804_ registers\[22\]\[53\] _13124_ VGND VGND VPWR VPWR _13128_ sky130_fd_sc_hd__mux2_1
XANTENNA_637 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26574_ _11598_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23786_ _10016_ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__buf_6
XANTENNA_648 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ registers\[8\]\[9\] registers\[9\]\[9\] registers\[10\]\[9\] registers\[11\]\[9\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__mux4_1
XANTENNA_659 _05196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28313_ registers\[2\]\[35\] _10378_ _12539_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1024 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25525_ _11043_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__clkbuf_1
X_22737_ _07385_ _09375_ _09376_ _07395_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__a22o_1
X_29293_ _09699_ registers\[22\]\[20\] _13091_ VGND VGND VPWR VPWR _13092_ sky130_fd_sc_hd__mux2_1
XFILLER_241_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28244_ registers\[2\]\[2\] _10309_ _12506_ VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__mux2_1
XFILLER_38_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25456_ _10860_ registers\[50\]\[62\] _10936_ VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__mux2_1
X_22668_ registers\[44\]\[57\] registers\[45\]\[57\] registers\[46\]\[57\] registers\[47\]\[57\]
+ _09078_ _09079_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__mux4_1
XFILLER_142_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24407_ net48 VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__buf_4
XFILLER_199_1128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21619_ registers\[44\]\[27\] registers\[45\]\[27\] registers\[46\]\[27\] registers\[47\]\[27\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__mux4_1
X_28175_ _12472_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__clkbuf_1
X_25387_ _10791_ registers\[50\]\[29\] _10959_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__mux2_1
X_22599_ registers\[28\]\[54\] registers\[29\]\[54\] registers\[30\]\[54\] registers\[31\]\[54\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__mux4_1
XFILLER_187_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27126_ _11919_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24338_ net24 VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__buf_4
XFILLER_193_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27057_ _11883_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24269_ _10320_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
X_26008_ _11299_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_218_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1003 _11832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_218_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1025 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18830_ registers\[44\]\[13\] registers\[45\]\[13\] registers\[46\]\[13\] registers\[47\]\[13\]
+ _05470_ _05471_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__mux4_1
XTAP_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1014 _12150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1025 _12647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1036 _13068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1047 _13281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1058 _13850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18761_ _05197_ _05511_ _05512_ _05202_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__a22o_1
XFILLER_62_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27959_ _12358_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__clkbuf_1
XTAP_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1069 _14347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ _14592_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__buf_6
XFILLER_23_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30970_ registers\[10\]\[47\] _13033_ _13966_ VGND VGND VPWR VPWR _13974_ sky130_fd_sc_hd__mux2_1
XFILLER_236_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ registers\[48\]\[9\] registers\[49\]\[9\] registers\[50\]\[9\] registers\[51\]\[9\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__mux4_1
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29629_ _13268_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__clkbuf_1
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17643_ registers\[24\]\[44\] registers\[25\]\[44\] registers\[26\]\[44\] registers\[27\]\[44\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__mux4_1
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32640_ clknet_leaf_267_CLK _00754_ VGND VGND VPWR VPWR registers\[58\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_17574_ _04355_ _04358_ _15974_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19313_ _06046_ _06049_ _05851_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__o21ba_1
X_16525_ _15003_ _15010_ _15017_ _15026_ VGND VGND VPWR VPWR _15027_ sky130_fd_sc_hd__or4_1
XFILLER_95_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32571_ clknet_leaf_305_CLK _00685_ VGND VGND VPWR VPWR registers\[5\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34310_ clknet_leaf_247_CLK _02424_ VGND VGND VPWR VPWR registers\[32\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31522_ _14264_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19244_ _05957_ _05966_ _05973_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__or4_4
X_16456_ _14951_ _14958_ _14959_ VGND VGND VPWR VPWR _14960_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35290_ clknet_leaf_7_CLK _03404_ VGND VGND VPWR VPWR registers\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34241_ clknet_leaf_257_CLK _02355_ VGND VGND VPWR VPWR registers\[33\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_31453_ _14205_ VGND VGND VPWR VPWR _14228_ sky130_fd_sc_hd__buf_4
X_19175_ registers\[20\]\[22\] registers\[21\]\[22\] registers\[22\]\[22\] registers\[23\]\[22\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__mux4_1
X_16387_ registers\[44\]\[9\] registers\[45\]\[9\] registers\[46\]\[9\] registers\[47\]\[9\]
+ _14512_ _14513_ VGND VGND VPWR VPWR _14892_ sky130_fd_sc_hd__mux4_1
XFILLER_247_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18126_ registers\[32\]\[59\] registers\[33\]\[59\] registers\[34\]\[59\] registers\[35\]\[59\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__mux4_1
XFILLER_160_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30404_ _13676_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__clkbuf_1
X_34172_ clknet_leaf_276_CLK _02286_ VGND VGND VPWR VPWR registers\[34\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31384_ registers\[7\]\[51\] net47 _14190_ VGND VGND VPWR VPWR _14192_ sky130_fd_sc_hd__mux2_1
XFILLER_157_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18057_ registers\[16\]\[56\] registers\[17\]\[56\] registers\[18\]\[56\] registers\[19\]\[56\]
+ _14602_ _14604_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__mux4_1
X_30335_ _13640_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__clkbuf_1
X_33123_ clknet_leaf_47_CLK _01237_ VGND VGND VPWR VPWR registers\[50\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17008_ registers\[16\]\[26\] registers\[17\]\[26\] registers\[18\]\[26\] registers\[19\]\[26\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15496_ sky130_fd_sc_hd__mux4_1
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33054_ clknet_leaf_37_CLK _01168_ VGND VGND VPWR VPWR registers\[51\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30266_ _13603_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32005_ clknet_leaf_28_CLK _00178_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30197_ _13567_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_1218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18959_ _05501_ _05704_ _05705_ _05506_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__a22o_1
XANTENNA_1570 _12860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_227_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1581 _14276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1592 _14539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21970_ registers\[32\]\[37\] registers\[33\]\[37\] registers\[34\]\[37\] registers\[35\]\[37\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__mux4_1
X_33956_ clknet_leaf_440_CLK _02070_ VGND VGND VPWR VPWR registers\[37\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32907_ clknet_leaf_166_CLK _01021_ VGND VGND VPWR VPWR registers\[54\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_20921_ _07313_ _07611_ _07612_ _07322_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__a22o_1
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33887_ clknet_leaf_16_CLK _02001_ VGND VGND VPWR VPWR registers\[38\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35626_ clknet_leaf_459_CLK _03740_ VGND VGND VPWR VPWR registers\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23640_ registers\[61\]\[36\] _09766_ _09976_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__mux2_1
X_32838_ clknet_leaf_194_CLK _00952_ VGND VGND VPWR VPWR registers\[55\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_20852_ _07325_ _07544_ _07545_ _07336_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__a22o_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23571_ registers\[61\]\[3\] _09664_ _09943_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__mux2_1
X_35557_ clknet_leaf_462_CLK _03671_ VGND VGND VPWR VPWR registers\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32769_ clknet_leaf_266_CLK _00883_ VGND VGND VPWR VPWR registers\[56\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_20783_ _07313_ _07477_ _07478_ _07322_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__a22o_1
XFILLER_23_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25310_ _10850_ registers\[51\]\[57\] _10920_ VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__mux2_1
X_22522_ registers\[0\]\[52\] registers\[1\]\[52\] registers\[2\]\[52\] registers\[3\]\[52\]
+ _09095_ _09096_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__mux4_1
X_34508_ clknet_leaf_148_CLK _02622_ VGND VGND VPWR VPWR registers\[2\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26290_ _11448_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35488_ clknet_leaf_468_CLK _03602_ VGND VGND VPWR VPWR registers\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_25241_ _10781_ registers\[51\]\[24\] _10887_ VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__mux2_1
X_22453_ _07369_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__buf_2
X_34439_ clknet_leaf_206_CLK _02553_ VGND VGND VPWR VPWR registers\[30\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_210_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_241_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21404_ _07392_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25172_ _10852_ registers\[52\]\[58\] _10836_ VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__mux2_1
XFILLER_157_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22384_ _09029_ _09034_ _08759_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__o21ba_1
XFILLER_163_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36109_ clknet_leaf_170_CLK _04223_ VGND VGND VPWR VPWR registers\[59\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_24123_ _09527_ registers\[58\]\[6\] _10233_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__mux2_1
XFILLER_135_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21335_ registers\[40\]\[19\] registers\[41\]\[19\] registers\[42\]\[19\] registers\[43\]\[19\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__mux4_1
XFILLER_203_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29980_ registers\[17\]\[26\] _12989_ _13446_ VGND VGND VPWR VPWR _13453_ sky130_fd_sc_hd__mux2_1
XFILLER_237_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28931_ registers\[24\]\[8\] _10321_ _12861_ VGND VGND VPWR VPWR _12870_ sky130_fd_sc_hd__mux2_1
X_24054_ _09594_ registers\[5\]\[38\] _10194_ VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__mux2_1
XFILLER_172_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21266_ registers\[44\]\[17\] registers\[45\]\[17\] registers\[46\]\[17\] registers\[47\]\[17\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__mux4_1
XFILLER_173_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_941 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23005_ _09598_ registers\[62\]\[40\] _09599_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__mux2_1
XFILLER_235_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20217_ registers\[60\]\[52\] registers\[61\]\[52\] registers\[62\]\[52\] registers\[63\]\[52\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28862_ _12833_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__clkbuf_1
X_21197_ registers\[36\]\[15\] registers\[37\]\[15\] registers\[38\]\[15\] registers\[39\]\[15\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__mux4_1
XFILLER_104_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20148_ registers\[0\]\[50\] registers\[1\]\[50\] registers\[2\]\[50\] registers\[3\]\[50\]
+ _06859_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__mux4_1
X_27813_ registers\[33\]\[54\] _10418_ _12277_ VGND VGND VPWR VPWR _12282_ sky130_fd_sc_hd__mux2_1
X_28793_ _12797_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__clkbuf_1
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20079_ registers\[12\]\[48\] registers\[13\]\[48\] registers\[14\]\[48\] registers\[15\]\[48\]
+ _06623_ _06624_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__mux4_1
X_24956_ _09615_ registers\[53\]\[48\] _10702_ VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__mux2_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27744_ registers\[33\]\[21\] _10349_ _12244_ VGND VGND VPWR VPWR _12246_ sky130_fd_sc_hd__mux2_1
XFILLER_218_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23907_ _10125_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
X_27675_ _12209_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_218_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24887_ _09546_ registers\[53\]\[15\] _10669_ VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__mux2_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_401 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29414_ _13155_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__clkbuf_1
X_26626_ _11625_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _10088_ VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__buf_4
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_434 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_445 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_456 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_467 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26557_ _11589_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__clkbuf_1
X_29345_ _09786_ registers\[22\]\[45\] _13113_ VGND VGND VPWR VPWR _13119_ sky130_fd_sc_hd__mux2_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23769_ _10052_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_478 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_489 _00165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16310_ registers\[40\]\[7\] registers\[41\]\[7\] registers\[42\]\[7\] registers\[43\]\[7\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14817_ sky130_fd_sc_hd__mux4_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25508_ registers\[4\]\[20\] _10346_ _11034_ VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__mux2_1
XFILLER_242_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29276_ _09683_ registers\[22\]\[12\] _13080_ VGND VGND VPWR VPWR _13083_ sky130_fd_sc_hd__mux2_1
X_17290_ registers\[24\]\[34\] registers\[25\]\[34\] registers\[26\]\[34\] registers\[27\]\[34\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15770_ sky130_fd_sc_hd__mux4_1
XFILLER_14_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26488_ _11552_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__clkbuf_1
X_16241_ registers\[32\]\[5\] registers\[33\]\[5\] registers\[34\]\[5\] registers\[35\]\[5\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14750_ sky130_fd_sc_hd__mux4_1
X_28227_ _12499_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__clkbuf_1
X_25439_ _10996_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16172_ _14660_ _14667_ _14674_ _14683_ VGND VGND VPWR VPWR _14684_ sky130_fd_sc_hd__or4_2
X_28158_ _12463_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_220_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27109_ _11816_ registers\[38\]\[41\] _11909_ VGND VGND VPWR VPWR _11911_ sky130_fd_sc_hd__mux2_1
X_28089_ _11849_ registers\[31\]\[57\] _12419_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__mux2_1
XFILLER_154_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30120_ _13526_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19931_ registers\[52\]\[44\] registers\[53\]\[44\] registers\[54\]\[44\] registers\[55\]\[44\]
+ _06369_ _06370_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__mux4_1
XFILLER_123_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30051_ registers\[17\]\[60\] _13060_ _13423_ VGND VGND VPWR VPWR _13490_ sky130_fd_sc_hd__mux2_1
X_19862_ registers\[48\]\[42\] registers\[49\]\[42\] registers\[50\]\[42\] registers\[51\]\[42\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__mux4_1
XFILLER_214_1117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput92 net92 VGND VGND VPWR VPWR D1[11] sky130_fd_sc_hd__buf_2
X_18813_ registers\[4\]\[12\] registers\[5\]\[12\] registers\[6\]\[12\] registers\[7\]\[12\]
+ _05423_ _05424_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__mux4_1
XFILLER_95_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19793_ _05120_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__buf_4
XTAP_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33810_ clknet_leaf_105_CLK _01924_ VGND VGND VPWR VPWR registers\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_18744_ registers\[24\]\[10\] registers\[25\]\[10\] registers\[26\]\[10\] registers\[27\]\[10\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__mux4_1
XTAP_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34790_ clknet_leaf_451_CLK _02904_ VGND VGND VPWR VPWR registers\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33741_ clknet_leaf_75_CLK _01855_ VGND VGND VPWR VPWR registers\[41\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_18675_ _05137_ _05428_ _05429_ _05147_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__a22o_1
X_30953_ registers\[10\]\[39\] _13016_ _13955_ VGND VGND VPWR VPWR _13965_ sky130_fd_sc_hd__mux2_1
XFILLER_237_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17626_ registers\[56\]\[44\] registers\[57\]\[44\] registers\[58\]\[44\] registers\[59\]\[44\]
+ _04408_ _15885_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__mux4_1
X_33672_ clknet_leaf_243_CLK _01786_ VGND VGND VPWR VPWR registers\[42\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30884_ registers\[10\]\[6\] _12947_ _13922_ VGND VGND VPWR VPWR _13929_ sky130_fd_sc_hd__mux2_1
XFILLER_17_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35411_ clknet_leaf_77_CLK _03525_ VGND VGND VPWR VPWR registers\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32623_ clknet_leaf_367_CLK _00737_ VGND VGND VPWR VPWR registers\[58\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17557_ registers\[36\]\[42\] registers\[37\]\[42\] registers\[38\]\[42\] registers\[39\]\[42\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__mux4_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_990 _11729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35342_ clknet_leaf_137_CLK _03456_ VGND VGND VPWR VPWR registers\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_16508_ _15006_ _15009_ _14934_ _14935_ VGND VGND VPWR VPWR _15010_ sky130_fd_sc_hd__o211a_2
XFILLER_147_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32554_ clknet_leaf_402_CLK _00668_ VGND VGND VPWR VPWR registers\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_17488_ _15892_ _15960_ _15961_ _15896_ VGND VGND VPWR VPWR _15962_ sky130_fd_sc_hd__a22o_1
XFILLER_220_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31505_ _14255_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__clkbuf_1
X_19227_ _05961_ _05965_ _05826_ _05827_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__o211a_1
X_35273_ clknet_leaf_155_CLK _03387_ VGND VGND VPWR VPWR registers\[17\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_16439_ registers\[4\]\[10\] registers\[5\]\[10\] registers\[6\]\[10\] registers\[7\]\[10\]
+ _14874_ _14875_ VGND VGND VPWR VPWR _14943_ sky130_fd_sc_hd__mux4_1
XFILLER_34_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32485_ clknet_leaf_450_CLK _00599_ VGND VGND VPWR VPWR registers\[60\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34224_ clknet_leaf_349_CLK _02338_ VGND VGND VPWR VPWR registers\[33\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_31436_ _14219_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__clkbuf_1
X_19158_ registers\[60\]\[22\] registers\[61\]\[22\] registers\[62\]\[22\] registers\[63\]\[22\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__mux4_1
XFILLER_191_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18109_ registers\[8\]\[58\] registers\[9\]\[58\] registers\[10\]\[58\] registers\[11\]\[58\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__mux4_1
X_31367_ registers\[7\]\[43\] net38 _14179_ VGND VGND VPWR VPWR _14183_ sky130_fd_sc_hd__mux2_1
X_34155_ clknet_leaf_425_CLK _02269_ VGND VGND VPWR VPWR registers\[34\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19089_ registers\[0\]\[20\] registers\[1\]\[20\] registers\[2\]\[20\] registers\[3\]\[20\]
+ _05830_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__mux4_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30318_ _13630_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__clkbuf_1
X_33106_ clknet_leaf_73_CLK _01220_ VGND VGND VPWR VPWR registers\[50\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_21120_ _07388_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__buf_4
XFILLER_105_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31298_ registers\[7\]\[10\] net2 _14146_ VGND VGND VPWR VPWR _14147_ sky130_fd_sc_hd__mux2_1
X_34086_ clknet_leaf_432_CLK _02200_ VGND VGND VPWR VPWR registers\[35\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_21051_ _07392_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__buf_4
X_33037_ clknet_leaf_140_CLK _01151_ VGND VGND VPWR VPWR registers\[52\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_30249_ _13594_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20002_ registers\[0\]\[46\] registers\[1\]\[46\] registers\[2\]\[46\] registers\[3\]\[46\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__mux4_1
XFILLER_119_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1075 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1048 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24810_ _10634_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25790_ _11185_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
X_34988_ clknet_leaf_403_CLK _03102_ VGND VGND VPWR VPWR registers\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_228_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_875 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24741_ _10586_ VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__buf_6
X_33939_ clknet_leaf_126_CLK _02053_ VGND VGND VPWR VPWR registers\[37\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21953_ registers\[12\]\[36\] registers\[13\]\[36\] registers\[14\]\[36\] registers\[15\]\[36\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__mux4_1
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_228_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ registers\[28\]\[6\] registers\[29\]\[6\] registers\[30\]\[6\] registers\[31\]\[6\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__mux4_1
X_27460_ _12095_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__clkbuf_1
X_24672_ _09603_ registers\[55\]\[42\] _10558_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__mux2_1
X_21884_ registers\[12\]\[34\] registers\[13\]\[34\] registers\[14\]\[34\] registers\[15\]\[34\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__mux4_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26411_ _11511_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ registers\[61\]\[28\] _09749_ _09965_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__mux2_1
X_35609_ clknet_leaf_14_CLK _03723_ VGND VGND VPWR VPWR registers\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_20835_ registers\[20\]\[4\] registers\[21\]\[4\] registers\[22\]\[4\] registers\[23\]\[4\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__mux4_1
X_27391_ registers\[36\]\[47\] _10403_ _12051_ VGND VGND VPWR VPWR _12059_ sky130_fd_sc_hd__mux2_1
XFILLER_70_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_247_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29130_ registers\[23\]\[25\] _12987_ _12977_ VGND VGND VPWR VPWR _12988_ sky130_fd_sc_hd__mux2_1
XFILLER_168_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26342_ _11475_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23554_ _09936_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20766_ _07377_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__buf_6
XFILLER_39_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22505_ registers\[32\]\[52\] registers\[33\]\[52\] registers\[34\]\[52\] registers\[35\]\[52\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__mux4_1
X_29061_ net34 VGND VGND VPWR VPWR _12941_ sky130_fd_sc_hd__buf_2
X_26273_ _10858_ registers\[44\]\[61\] _11371_ VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__mux2_1
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23485_ _09900_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
X_20697_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__buf_4
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28012_ _11771_ registers\[31\]\[20\] _12386_ VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25224_ _10764_ registers\[51\]\[16\] _10876_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__mux2_1
X_22436_ registers\[56\]\[50\] registers\[57\]\[50\] registers\[58\]\[50\] registers\[59\]\[50\]
+ _08880_ _09013_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__mux4_1
XFILLER_202_1054 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25155_ _10841_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22367_ _07284_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_191_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_191_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_100_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24106_ _09646_ registers\[5\]\[63\] _10160_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__mux2_1
XFILLER_184_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21318_ registers\[0\]\[18\] registers\[1\]\[18\] registers\[2\]\[18\] registers\[3\]\[18\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__mux4_1
XFILLER_174_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25086_ _10793_ registers\[52\]\[30\] _10794_ VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__mux2_1
X_29963_ registers\[17\]\[18\] _12972_ _13435_ VGND VGND VPWR VPWR _13444_ sky130_fd_sc_hd__mux2_1
XFILLER_190_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22298_ _08677_ _08947_ _08950_ _08681_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__a22o_1
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28914_ _12860_ VGND VGND VPWR VPWR _12861_ sky130_fd_sc_hd__buf_4
XFILLER_2_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24037_ _10160_ VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__buf_6
XFILLER_215_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21249_ _07366_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29894_ _13407_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_996 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28845_ _11795_ registers\[25\]\[31\] _12823_ VGND VGND VPWR VPWR _12825_ sky130_fd_sc_hd__mux2_1
XFILLER_93_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16790_ _15139_ _15280_ _15283_ _15142_ VGND VGND VPWR VPWR _15284_ sky130_fd_sc_hd__a22o_1
X_28776_ _11861_ registers\[26\]\[63\] _12718_ VGND VGND VPWR VPWR _12788_ sky130_fd_sc_hd__mux2_1
X_25988_ _11289_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_246_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24939_ _10657_ VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__buf_4
X_27727_ registers\[33\]\[13\] _10332_ _12233_ VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__mux2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18460_ registers\[4\]\[2\] registers\[5\]\[2\] registers\[6\]\[2\] registers\[7\]\[2\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux4_1
XFILLER_2_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27658_ _12200_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_220 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _14541_ VGND VGND VPWR VPWR _15887_ sky130_fd_sc_hd__buf_4
XFILLER_233_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_253 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18391_ registers\[28\]\[0\] registers\[29\]\[0\] registers\[30\]\[0\] registers\[31\]\[0\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__mux4_1
X_26609_ _11616_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__clkbuf_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27589_ _12164_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_264 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_286 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _14546_ VGND VGND VPWR VPWR _15820_ sky130_fd_sc_hd__clkbuf_8
XFILLER_158_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_297 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29328_ _09769_ registers\[22\]\[37\] _13102_ VGND VGND VPWR VPWR _13110_ sky130_fd_sc_hd__mux2_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17273_ registers\[56\]\[34\] registers\[57\]\[34\] registers\[58\]\[34\] registers\[59\]\[34\]
+ _15752_ _15542_ VGND VGND VPWR VPWR _15753_ sky130_fd_sc_hd__mux4_1
X_29259_ _09666_ registers\[22\]\[4\] _13069_ VGND VGND VPWR VPWR _13074_ sky130_fd_sc_hd__mux2_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16224_ _14558_ _14732_ _14733_ _14568_ VGND VGND VPWR VPWR _14734_ sky130_fd_sc_hd__a22o_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19012_ registers\[60\]\[18\] registers\[61\]\[18\] registers\[62\]\[18\] registers\[63\]\[18\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__mux4_1
X_32270_ clknet_leaf_113_CLK _00384_ VGND VGND VPWR VPWR registers\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31221_ registers\[8\]\[38\] net32 _14097_ VGND VGND VPWR VPWR _14106_ sky130_fd_sc_hd__mux2_1
X_16155_ _14663_ _14666_ _14554_ _14556_ VGND VGND VPWR VPWR _14667_ sky130_fd_sc_hd__o211a_1
XFILLER_31_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_182_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_182_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31152_ registers\[8\]\[5\] net56 _14064_ VGND VGND VPWR VPWR _14070_ sky130_fd_sc_hd__mux2_1
X_16086_ _14509_ VGND VGND VPWR VPWR _14600_ sky130_fd_sc_hd__buf_12
XFILLER_6_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30103_ registers\[16\]\[20\] _12976_ _13517_ VGND VGND VPWR VPWR _13518_ sky130_fd_sc_hd__mux2_1
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19914_ _06530_ _06632_ _06633_ _06535_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__a22o_1
XFILLER_29_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35960_ clknet_leaf_314_CLK _04074_ VGND VGND VPWR VPWR registers\[6\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_31083_ _14033_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30034_ _13481_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__clkbuf_1
X_34911_ clknet_leaf_488_CLK _03025_ VGND VGND VPWR VPWR registers\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19845_ _06563_ _06566_ _06537_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__o21ba_1
XFILLER_122_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35891_ clknet_leaf_380_CLK _04005_ VGND VGND VPWR VPWR registers\[7\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34842_ clknet_leaf_0_CLK _02956_ VGND VGND VPWR VPWR registers\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_19776_ _05095_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__buf_4
XFILLER_56_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16988_ registers\[60\]\[26\] registers\[61\]\[26\] registers\[62\]\[26\] registers\[63\]\[26\]
+ _15413_ _15207_ VGND VGND VPWR VPWR _15476_ sky130_fd_sc_hd__mux4_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18727_ registers\[60\]\[10\] registers\[61\]\[10\] registers\[62\]\[10\] registers\[63\]\[10\]
+ _05276_ _05413_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__mux4_1
XFILLER_225_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34773_ clknet_leaf_88_CLK _02887_ VGND VGND VPWR VPWR registers\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31985_ clknet_leaf_22_CLK _00156_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
X_33724_ clknet_leaf_277_CLK _01838_ VGND VGND VPWR VPWR registers\[41\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_236_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18658_ _05092_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__buf_4
X_30936_ _13956_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1087 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17609_ registers\[24\]\[43\] registers\[25\]\[43\] registers\[26\]\[43\] registers\[27\]\[43\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__mux4_1
XFILLER_24_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33655_ clknet_leaf_341_CLK _01769_ VGND VGND VPWR VPWR registers\[42\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_30867_ _13919_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__clkbuf_1
X_18589_ registers\[8\]\[6\] registers\[9\]\[6\] registers\[10\]\[6\] registers\[11\]\[6\]
+ _05312_ _05313_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__mux4_1
XFILLER_36_1303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20620_ _07278_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__buf_4
X_32606_ clknet_leaf_38_CLK _00720_ VGND VGND VPWR VPWR registers\[58\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33586_ clknet_leaf_361_CLK _01700_ VGND VGND VPWR VPWR registers\[43\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_30798_ _13883_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_966 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35325_ clknet_leaf_179_CLK _03439_ VGND VGND VPWR VPWR registers\[16\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20551_ _07247_ _07250_ _05073_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__o21ba_1
XFILLER_123_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32537_ clknet_leaf_475_CLK _00651_ VGND VGND VPWR VPWR registers\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35256_ clknet_leaf_428_CLK _03370_ VGND VGND VPWR VPWR registers\[17\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_23270_ net35 VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__buf_4
X_20482_ _07181_ _07184_ _05162_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__o21ba_1
XFILLER_192_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32468_ clknet_leaf_63_CLK _00582_ VGND VGND VPWR VPWR registers\[60\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22221_ registers\[44\]\[44\] registers\[45\]\[44\] registers\[46\]\[44\] registers\[47\]\[44\]
+ _08735_ _08736_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__mux4_1
X_34207_ clknet_leaf_16_CLK _02321_ VGND VGND VPWR VPWR registers\[33\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_31419_ _14210_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_173_CLK clknet_6_25__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_173_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35187_ clknet_leaf_421_CLK _03301_ VGND VGND VPWR VPWR registers\[18\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_32399_ clknet_leaf_110_CLK _00513_ VGND VGND VPWR VPWR registers\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1085 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22152_ registers\[32\]\[42\] registers\[33\]\[42\] registers\[34\]\[42\] registers\[35\]\[42\]
+ _08702_ _08703_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__mux4_1
X_34138_ clknet_leaf_18_CLK _02252_ VGND VGND VPWR VPWR registers\[34\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21103_ registers\[48\]\[12\] registers\[49\]\[12\] registers\[50\]\[12\] registers\[51\]\[12\]
+ _07643_ _07644_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__mux4_1
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34069_ clknet_leaf_121_CLK _02183_ VGND VGND VPWR VPWR registers\[35\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_26960_ _11822_ registers\[3\]\[44\] _11814_ VGND VGND VPWR VPWR _11823_ sky130_fd_sc_hd__mux2_1
X_22083_ registers\[56\]\[40\] registers\[57\]\[40\] registers\[58\]\[40\] registers\[59\]\[40\]
+ _08537_ _08670_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__mux4_1
XTAP_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25911_ _10766_ registers\[46\]\[17\] _11241_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__mux2_1
X_21034_ _07347_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__buf_6
X_26891_ net15 VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__clkbuf_4
XFILLER_219_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28630_ _12711_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__clkbuf_1
X_25842_ _11212_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_44__f_CLK clknet_5_22_0_CLK VGND VGND VPWR VPWR clknet_6_44__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25773_ _11176_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
X_28561_ _12675_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__clkbuf_1
X_22985_ net28 VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24724_ _10589_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
X_27512_ _11813_ registers\[35\]\[40\] _12122_ VGND VGND VPWR VPWR _12123_ sky130_fd_sc_hd__mux2_1
X_28492_ _11847_ registers\[28\]\[56\] _12632_ VGND VGND VPWR VPWR _12639_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21936_ _08469_ _08597_ _08598_ _08472_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__a22o_1
XFILLER_103_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27443_ _12086_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24655_ _09586_ registers\[55\]\[34\] _10547_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__mux2_1
XFILLER_231_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21867_ _08462_ _08530_ _08531_ _08467_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__a22o_1
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_231_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _09942_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__buf_4
X_20818_ registers\[60\]\[4\] registers\[61\]\[4\] registers\[62\]\[4\] registers\[63\]\[4\]
+ _07512_ _07329_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__mux4_1
X_27374_ registers\[36\]\[39\] _10386_ _12040_ VGND VGND VPWR VPWR _12050_ sky130_fd_sc_hd__mux2_1
X_24586_ _09517_ registers\[55\]\[1\] _10514_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__mux2_1
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21798_ registers\[40\]\[32\] registers\[41\]\[32\] registers\[42\]\[32\] registers\[43\]\[32\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__mux4_1
X_29113_ net13 VGND VGND VPWR VPWR _12976_ sky130_fd_sc_hd__clkbuf_4
X_26325_ _10775_ registers\[43\]\[21\] _11465_ VGND VGND VPWR VPWR _11467_ sky130_fd_sc_hd__mux2_1
X_23537_ _09624_ registers\[19\]\[52\] _09925_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__mux2_1
XFILLER_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20749_ registers\[56\]\[2\] registers\[57\]\[2\] registers\[58\]\[2\] registers\[59\]\[2\]
+ _07315_ _07317_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__mux4_1
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29044_ registers\[24\]\[62\] _10434_ _12860_ VGND VGND VPWR VPWR _12929_ sky130_fd_sc_hd__mux2_1
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26256_ _11430_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
X_23468_ _09891_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25207_ _10747_ registers\[51\]\[8\] _10865_ VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__mux2_1
X_22419_ _08761_ _09067_ _09068_ _08764_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__a22o_1
XFILLER_13_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_164_CLK clknet_6_30__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_164_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26187_ _11371_ VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__buf_4
X_23399_ registers\[39\]\[52\] _09802_ _09851_ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__mux2_1
XFILLER_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25138_ _10829_ registers\[52\]\[47\] _10815_ VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__mux2_1
XFILLER_100_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17960_ _04486_ _04732_ _04733_ _04489_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__a22o_1
XFILLER_139_1379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29946_ _13423_ VGND VGND VPWR VPWR _13435_ sky130_fd_sc_hd__buf_4
X_25069_ net18 VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__buf_2
XFILLER_151_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16911_ _15401_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
X_17891_ _04663_ _04666_ _04630_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__o21ba_1
X_29877_ registers\[18\]\[41\] _13021_ _13397_ VGND VGND VPWR VPWR _13399_ sky130_fd_sc_hd__mux2_1
XFILLER_215_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19630_ _06357_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__buf_2
XFILLER_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28828_ _11778_ registers\[25\]\[23\] _12812_ VGND VGND VPWR VPWR _12816_ sky130_fd_sc_hd__mux2_1
X_16842_ _14527_ VGND VGND VPWR VPWR _15334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_120_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19561_ _06187_ _06289_ _06290_ _06192_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a22o_1
X_28759_ _12779_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__clkbuf_1
X_16773_ registers\[36\]\[20\] registers\[37\]\[20\] registers\[38\]\[20\] registers\[39\]\[20\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15267_ sky130_fd_sc_hd__mux4_1
XFILLER_46_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18512_ _05267_ _05270_ _05074_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31770_ registers\[59\]\[42\] net37 _14392_ VGND VGND VPWR VPWR _14395_ sky130_fd_sc_hd__mux2_1
X_19492_ _06220_ _06223_ _06194_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__o21ba_1
XFILLER_92_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30721_ registers\[12\]\[57\] _13054_ _13835_ VGND VGND VPWR VPWR _13843_ sky130_fd_sc_hd__mux2_1
X_18443_ _05059_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__buf_6
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33440_ clknet_leaf_34_CLK _01554_ VGND VGND VPWR VPWR registers\[45\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_18374_ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__buf_4
X_30652_ registers\[12\]\[24\] _12985_ _13802_ VGND VGND VPWR VPWR _13807_ sky130_fd_sc_hd__mux2_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17325_ registers\[28\]\[35\] registers\[29\]\[35\] registers\[30\]\[35\] registers\[31\]\[35\]
+ _15707_ _15708_ VGND VGND VPWR VPWR _15804_ sky130_fd_sc_hd__mux4_1
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30583_ _13770_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__clkbuf_1
X_33371_ clknet_leaf_30_CLK _01485_ VGND VGND VPWR VPWR registers\[46\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35110_ clknet_leaf_463_CLK _03224_ VGND VGND VPWR VPWR registers\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_32322_ clknet_leaf_222_CLK _00436_ VGND VGND VPWR VPWR registers\[19\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36090_ clknet_leaf_284_CLK _04204_ VGND VGND VPWR VPWR registers\[59\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_17256_ registers\[24\]\[33\] registers\[25\]\[33\] registers\[26\]\[33\] registers\[27\]\[33\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15737_ sky130_fd_sc_hd__mux4_1
XFILLER_146_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16207_ registers\[32\]\[4\] registers\[33\]\[4\] registers\[34\]\[4\] registers\[35\]\[4\]
+ _14519_ _14521_ VGND VGND VPWR VPWR _14717_ sky130_fd_sc_hd__mux4_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35041_ clknet_leaf_489_CLK _03155_ VGND VGND VPWR VPWR registers\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_155_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_155_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32253_ clknet_leaf_268_CLK _00367_ VGND VGND VPWR VPWR registers\[39\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_17187_ registers\[16\]\[31\] registers\[17\]\[31\] registers\[18\]\[31\] registers\[19\]\[31\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15670_ sky130_fd_sc_hd__mux4_1
XFILLER_143_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16138_ _14496_ VGND VGND VPWR VPWR _14650_ sky130_fd_sc_hd__buf_6
X_31204_ _14063_ VGND VGND VPWR VPWR _14097_ sky130_fd_sc_hd__buf_4
X_32184_ clknet_leaf_485_CLK _00298_ VGND VGND VPWR VPWR registers\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31135_ _14060_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__clkbuf_1
X_16069_ _14570_ _14575_ _14580_ _14582_ VGND VGND VPWR VPWR _14583_ sky130_fd_sc_hd__a22o_1
XFILLER_170_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35943_ clknet_leaf_457_CLK _04057_ VGND VGND VPWR VPWR registers\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_31066_ _14024_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30017_ _13472_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19828_ registers\[60\]\[41\] registers\[61\]\[41\] registers\[62\]\[41\] registers\[63\]\[41\]
+ _06305_ _06442_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__mux4_1
XFILLER_111_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35874_ clknet_leaf_469_CLK _03988_ VGND VGND VPWR VPWR registers\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34825_ clknet_leaf_220_CLK _02939_ VGND VGND VPWR VPWR registers\[24\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19759_ _06374_ _06481_ _06482_ _06377_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__a22o_1
XFILLER_216_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34756_ clknet_leaf_219_CLK _02870_ VGND VGND VPWR VPWR registers\[25\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_22770_ registers\[0\]\[60\] registers\[1\]\[60\] registers\[2\]\[60\] registers\[3\]\[60\]
+ _07406_ _07407_ VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__mux4_1
XFILLER_209_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31968_ clknet_leaf_4_CLK _00137_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_1
XFILLER_224_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21721_ registers\[32\]\[30\] registers\[33\]\[30\] registers\[34\]\[30\] registers\[35\]\[30\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__mux4_1
X_33707_ clknet_leaf_428_CLK _01821_ VGND VGND VPWR VPWR registers\[41\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30919_ _13947_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__clkbuf_1
X_34687_ clknet_leaf_189_CLK _02801_ VGND VGND VPWR VPWR registers\[26\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31899_ _14462_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__clkbuf_1
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24440_ net60 VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__clkbuf_4
XFILLER_244_1441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33638_ clknet_leaf_57_CLK _01752_ VGND VGND VPWR VPWR registers\[42\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_21652_ registers\[36\]\[28\] registers\[37\]\[28\] registers\[38\]\[28\] registers\[39\]\[28\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__mux4_1
XFILLER_71_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _07301_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__buf_4
XFILLER_21_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24371_ registers\[57\]\[40\] _10388_ _10389_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__mux2_1
XFILLER_178_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_394_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_394_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21583_ _08126_ _08254_ _08255_ _08129_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__a22o_1
X_33569_ clknet_leaf_39_CLK _01683_ VGND VGND VPWR VPWR registers\[43\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26110_ _11353_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
X_23322_ net52 VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__buf_4
X_35308_ clknet_leaf_396_CLK _03422_ VGND VGND VPWR VPWR registers\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_20534_ _05060_ _07233_ _07234_ _05066_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__a22o_1
XFILLER_220_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27090_ _11797_ registers\[38\]\[32\] _11898_ VGND VGND VPWR VPWR _11901_ sky130_fd_sc_hd__mux2_1
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26041_ _11317_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23253_ net29 VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__clkbuf_4
X_35239_ clknet_leaf_448_CLK _03353_ VGND VGND VPWR VPWR registers\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_146_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_146_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20465_ registers\[60\]\[60\] registers\[61\]\[60\] registers\[62\]\[60\] registers\[63\]\[60\]
+ _06991_ _05143_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__mux4_1
XFILLER_134_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_229_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22204_ _07305_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__buf_4
XFILLER_165_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23184_ _09708_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__buf_4
X_20396_ registers\[32\]\[58\] registers\[33\]\[58\] registers\[34\]\[58\] registers\[35\]\[58\]
+ _06809_ _06810_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__mux4_1
X_29800_ _13358_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__clkbuf_1
X_22135_ registers\[12\]\[41\] registers\[13\]\[41\] registers\[14\]\[41\] registers\[15\]\[41\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__mux4_1
XTAP_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput260 net260 VGND VGND VPWR VPWR D3[48] sky130_fd_sc_hd__buf_2
X_27992_ _12376_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__clkbuf_1
XTAP_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput271 net271 VGND VGND VPWR VPWR D3[58] sky130_fd_sc_hd__buf_2
XFILLER_245_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29731_ registers\[1\]\[36\] _13010_ _13315_ VGND VGND VPWR VPWR _13322_ sky130_fd_sc_hd__mux2_1
X_22066_ _08418_ _08724_ _08725_ _08421_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__a22o_1
X_26943_ net33 VGND VGND VPWR VPWR _11811_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21017_ _07287_ VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__buf_4
XTAP_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29662_ registers\[1\]\[3\] _12941_ _13282_ VGND VGND VPWR VPWR _13286_ sky130_fd_sc_hd__mux2_1
XFILLER_48_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26874_ _11764_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28613_ _12702_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25825_ _10814_ registers\[47\]\[40\] _11203_ VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__mux2_1
X_29593_ _13249_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_114_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25756_ _11167_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28544_ _12666_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__clkbuf_1
X_22968_ _09574_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_1216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24707_ _09638_ registers\[55\]\[59\] _10569_ VGND VGND VPWR VPWR _10579_ sky130_fd_sc_hd__mux2_1
X_21919_ registers\[4\]\[35\] registers\[5\]\[35\] registers\[6\]\[35\] registers\[7\]\[35\]
+ _08345_ _08346_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__mux4_1
XFILLER_215_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25687_ _11085_ VGND VGND VPWR VPWR _11130_ sky130_fd_sc_hd__buf_4
X_28475_ _11830_ registers\[28\]\[48\] _12621_ VGND VGND VPWR VPWR _12630_ sky130_fd_sc_hd__mux2_1
X_22899_ _09527_ registers\[62\]\[6\] _09515_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__mux2_1
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27426_ _11863_ _09868_ VGND VGND VPWR VPWR _12077_ sky130_fd_sc_hd__nand2_8
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24638_ _09569_ registers\[55\]\[26\] _10536_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__mux2_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_230_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_763 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24569_ _09638_ registers\[56\]\[59\] _10495_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_385_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_385_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27357_ _12041_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_212_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17110_ _15591_ _15594_ _15288_ VGND VGND VPWR VPWR _15595_ sky130_fd_sc_hd__o21ba_1
XFILLER_106_1356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_211_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18090_ registers\[20\]\[57\] registers\[21\]\[57\] registers\[22\]\[57\] registers\[23\]\[57\]
+ _04639_ _04640_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux4_1
XFILLER_129_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26308_ _10758_ registers\[43\]\[13\] _11454_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__mux2_1
X_27288_ _12004_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17041_ _15290_ _15526_ _15527_ _15293_ VGND VGND VPWR VPWR _15528_ sky130_fd_sc_hd__a22o_1
X_29027_ _12920_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26239_ _11421_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_137_CLK clknet_6_22__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_137_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18992_ _05734_ _05737_ _05508_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__o21ba_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ registers\[36\]\[53\] registers\[37\]\[53\] registers\[38\]\[53\] registers\[39\]\[53\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__mux4_1
X_29929_ _13426_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32940_ clknet_leaf_370_CLK _01054_ VGND VGND VPWR VPWR registers\[53\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17874_ registers\[44\]\[51\] registers\[45\]\[51\] registers\[46\]\[51\] registers\[47\]\[51\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__mux4_1
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19613_ _05051_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__clkbuf_8
XFILLER_120_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16825_ _15314_ _15317_ _15277_ _15278_ VGND VGND VPWR VPWR _15318_ sky130_fd_sc_hd__o211a_1
X_32871_ clknet_leaf_437_CLK _00985_ VGND VGND VPWR VPWR registers\[54\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34610_ clknet_leaf_409_CLK _02724_ VGND VGND VPWR VPWR registers\[27\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_31822_ _14422_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__clkbuf_1
X_19544_ registers\[52\]\[33\] registers\[53\]\[33\] registers\[54\]\[33\] registers\[55\]\[33\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__mux4_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35590_ clknet_leaf_211_CLK _03704_ VGND VGND VPWR VPWR registers\[12\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_16756_ _15144_ _15249_ _15250_ _15147_ VGND VGND VPWR VPWR _15251_ sky130_fd_sc_hd__a22o_1
XFILLER_228_1403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_222_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34541_ clknet_leaf_402_CLK _02655_ VGND VGND VPWR VPWR registers\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_31753_ registers\[59\]\[34\] net28 _14381_ VGND VGND VPWR VPWR _14386_ sky130_fd_sc_hd__mux2_1
X_19475_ registers\[60\]\[31\] registers\[61\]\[31\] registers\[62\]\[31\] registers\[63\]\[31\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__mux4_1
X_16687_ registers\[16\]\[17\] registers\[17\]\[17\] registers\[18\]\[17\] registers\[19\]\[17\]
+ _15151_ _15152_ VGND VGND VPWR VPWR _15184_ sky130_fd_sc_hd__mux4_1
X_18426_ _05184_ _05187_ _05134_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__o21ba_1
X_30704_ registers\[12\]\[49\] _13037_ _13824_ VGND VGND VPWR VPWR _13834_ sky130_fd_sc_hd__mux2_1
X_34472_ clknet_leaf_457_CLK _02586_ VGND VGND VPWR VPWR registers\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31684_ registers\[59\]\[1\] net12 _14348_ VGND VGND VPWR VPWR _14350_ sky130_fd_sc_hd__mux2_1
XFILLER_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_222_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36211_ clknet_leaf_115_CLK _00094_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dfxtp_1
X_33423_ clknet_leaf_131_CLK _01537_ VGND VGND VPWR VPWR registers\[45\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_221_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18357_ _05041_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__buf_12
X_30635_ registers\[12\]\[16\] _12968_ _13791_ VGND VGND VPWR VPWR _13798_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_376_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_376_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17308_ _15541_ _15785_ _15786_ _15547_ VGND VGND VPWR VPWR _15787_ sky130_fd_sc_hd__a22o_1
X_36142_ clknet_leaf_365_CLK _04256_ VGND VGND VPWR VPWR registers\[49\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_33354_ clknet_leaf_163_CLK _01468_ VGND VGND VPWR VPWR registers\[47\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18288_ _05041_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__buf_12
X_30566_ _13761_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_8__f_CLK clknet_5_4_0_CLK VGND VGND VPWR VPWR clknet_6_8__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32305_ clknet_leaf_396_CLK _00419_ VGND VGND VPWR VPWR registers\[19\]\[35\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_128_CLK clknet_6_23__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_128_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17239_ _15716_ _15719_ _15612_ VGND VGND VPWR VPWR _15720_ sky130_fd_sc_hd__o21ba_1
X_36073_ clknet_leaf_423_CLK _04187_ VGND VGND VPWR VPWR registers\[59\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_33285_ clknet_leaf_258_CLK _01399_ VGND VGND VPWR VPWR registers\[48\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30497_ _13725_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35024_ clknet_leaf_114_CLK _03138_ VGND VGND VPWR VPWR registers\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20250_ registers\[52\]\[53\] registers\[53\]\[53\] registers\[54\]\[53\] registers\[55\]\[53\]
+ _06712_ _06713_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__mux4_1
XFILLER_7_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32236_ clknet_leaf_379_CLK _00350_ VGND VGND VPWR VPWR registers\[39\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20181_ registers\[60\]\[51\] registers\[61\]\[51\] registers\[62\]\[51\] registers\[63\]\[51\]
+ _06648_ _06785_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__mux4_1
XFILLER_118_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32167_ clknet_leaf_108_CLK _00281_ VGND VGND VPWR VPWR registers\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31118_ registers\[0\]\[53\] _13046_ _14048_ VGND VGND VPWR VPWR _14052_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32098_ clknet_leaf_484_CLK _00012_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23940_ _10142_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_300_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_300_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35926_ clknet_leaf_83_CLK _04040_ VGND VGND VPWR VPWR registers\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_31049_ registers\[0\]\[20\] _12976_ _14015_ VGND VGND VPWR VPWR _14016_ sky130_fd_sc_hd__mux2_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35857_ clknet_leaf_76_CLK _03971_ VGND VGND VPWR VPWR registers\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23871_ _10106_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25610_ registers\[48\]\[3\] _10311_ _11086_ VGND VGND VPWR VPWR _11090_ sky130_fd_sc_hd__mux2_1
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22822_ registers\[56\]\[62\] registers\[57\]\[62\] registers\[58\]\[62\] registers\[59\]\[62\]
+ _09223_ _07388_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__mux4_1
X_34808_ clknet_leaf_314_CLK _02922_ VGND VGND VPWR VPWR registers\[24\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_26590_ _11606_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__clkbuf_1
X_35788_ clknet_leaf_149_CLK _03902_ VGND VGND VPWR VPWR registers\[0\]\[62\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_808 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_819 _09118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_25541_ registers\[4\]\[36\] _10380_ _11045_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__mux2_1
X_22753_ _09371_ _09378_ _09385_ _09392_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__or4_4
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34739_ clknet_leaf_409_CLK _02853_ VGND VGND VPWR VPWR registers\[25\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28260_ _12505_ VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__buf_4
X_21704_ registers\[8\]\[29\] registers\[9\]\[29\] registers\[10\]\[29\] registers\[11\]\[29\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__mux4_1
XFILLER_53_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25472_ registers\[4\]\[3\] _10311_ _11012_ VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__mux2_1
XFILLER_80_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22684_ _07296_ _09324_ _09325_ _07302_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__a22o_1
XFILLER_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24423_ registers\[57\]\[57\] _10424_ _10410_ VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__mux2_1
X_27211_ _11964_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__clkbuf_1
X_21635_ registers\[12\]\[27\] registers\[13\]\[27\] registers\[14\]\[27\] registers\[15\]\[27\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__mux4_1
X_28191_ _11816_ registers\[30\]\[41\] _12479_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__mux2_1
XFILLER_233_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_367_CLK clknet_6_42__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_367_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_240_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27142_ _11849_ registers\[38\]\[57\] _11920_ VGND VGND VPWR VPWR _11928_ sky130_fd_sc_hd__mux2_1
XFILLER_138_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24354_ net29 VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__buf_4
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21566_ registers\[4\]\[25\] registers\[5\]\[25\] registers\[6\]\[25\] registers\[7\]\[25\]
+ _08002_ _08003_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__mux4_1
XFILLER_165_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23305_ registers\[9\]\[50\] _09797_ _09798_ VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__mux2_1
XFILLER_193_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_119_CLK clknet_6_21__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_119_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20517_ _05077_ _07216_ _07217_ _05086_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a22o_1
XFILLER_165_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27073_ _11780_ registers\[38\]\[24\] _11887_ VGND VGND VPWR VPWR _11892_ sky130_fd_sc_hd__mux2_1
X_24285_ _10331_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21497_ _07303_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__buf_4
X_26024_ _11308_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23236_ _09752_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20448_ _06868_ _07150_ _07151_ _06871_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__a22o_1
XTAP_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_1275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_877 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23167_ registers\[9\]\[3\] _09664_ _09709_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__mux2_1
XFILLER_49_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20379_ registers\[8\]\[57\] registers\[9\]\[57\] registers\[10\]\[57\] registers\[11\]\[57\]
+ _05052_ _05054_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__mux4_1
XTAP_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1207 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22118_ registers\[40\]\[41\] registers\[41\]\[41\] registers\[42\]\[41\] registers\[43\]\[41\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__mux4_1
XTAP_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1218 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23098_ _09665_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__clkbuf_1
XTAP_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27975_ _12367_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1229 _00030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29714_ registers\[1\]\[28\] _12993_ _13304_ VGND VGND VPWR VPWR _13313_ sky130_fd_sc_hd__mux2_1
XTAP_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26926_ _11799_ registers\[3\]\[33\] _11793_ VGND VGND VPWR VPWR _11800_ sky130_fd_sc_hd__mux2_1
X_22049_ _08705_ _08708_ _08397_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__o21ba_1
XTAP_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29645_ _13276_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__clkbuf_1
XTAP_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26857_ net3 VGND VGND VPWR VPWR _11753_ sky130_fd_sc_hd__buf_4
XFILLER_36_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16610_ registers\[0\]\[15\] registers\[1\]\[15\] registers\[2\]\[15\] registers\[3\]\[15\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _15109_ sky130_fd_sc_hd__mux4_1
X_25808_ _10798_ registers\[47\]\[32\] _11192_ VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__mux2_1
XFILLER_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17590_ registers\[36\]\[43\] registers\[37\]\[43\] registers\[38\]\[43\] registers\[39\]\[43\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__mux4_1
X_29576_ _13240_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__clkbuf_1
X_26788_ registers\[40\]\[48\] _10405_ _11702_ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28527_ _12657_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16541_ registers\[8\]\[13\] registers\[9\]\[13\] registers\[10\]\[13\] registers\[11\]\[13\]
+ _14763_ _14764_ VGND VGND VPWR VPWR _15042_ sky130_fd_sc_hd__mux4_1
X_25739_ _10510_ _11157_ VGND VGND VPWR VPWR _11158_ sky130_fd_sc_hd__nand2_8
XFILLER_56_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19260_ _05051_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__buf_4
X_28458_ _12576_ VGND VGND VPWR VPWR _12621_ sky130_fd_sc_hd__clkbuf_8
X_16472_ _14971_ _14974_ _14934_ _14935_ VGND VGND VPWR VPWR _14975_ sky130_fd_sc_hd__o211a_2
XFILLER_143_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18211_ _14570_ _04975_ _04976_ _14582_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a22o_1
X_27409_ _12068_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_358_CLK clknet_6_43__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_358_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19191_ registers\[52\]\[23\] registers\[53\]\[23\] registers\[54\]\[23\] registers\[55\]\[23\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__mux4_1
X_28389_ _11744_ registers\[28\]\[7\] _12577_ VGND VGND VPWR VPWR _12585_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18142_ registers\[12\]\[59\] registers\[13\]\[59\] registers\[14\]\[59\] registers\[15\]\[59\]
+ _04730_ _04731_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__mux4_1
XFILLER_12_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30420_ _09780_ registers\[14\]\[42\] _13682_ VGND VGND VPWR VPWR _13685_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1017 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18073_ registers\[48\]\[57\] registers\[49\]\[57\] registers\[50\]\[57\] registers\[51\]\[57\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__mux4_1
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30351_ _13648_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17024_ _15505_ _15510_ _15269_ VGND VGND VPWR VPWR _15511_ sky130_fd_sc_hd__o21ba_1
X_33070_ clknet_leaf_365_CLK _01184_ VGND VGND VPWR VPWR registers\[51\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_30282_ registers\[15\]\[41\] _13021_ _13610_ VGND VGND VPWR VPWR _13612_ sky130_fd_sc_hd__mux2_1
XFILLER_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32021_ clknet_leaf_181_CLK _00199_ VGND VGND VPWR VPWR registers\[62\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ registers\[60\]\[17\] registers\[61\]\[17\] registers\[62\]\[17\] registers\[63\]\[17\]
+ _05619_ _05413_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__mux4_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1730 _00178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1741 _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17926_ _04486_ _04699_ _04700_ _04489_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__a22o_1
XANTENNA_1752 _06979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33972_ clknet_leaf_350_CLK _02086_ VGND VGND VPWR VPWR registers\[37\]\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1763 _07795_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1774 _11657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35711_ clknet_leaf_296_CLK _03825_ VGND VGND VPWR VPWR registers\[10\]\[49\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1785 _14518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32923_ clknet_leaf_57_CLK _01037_ VGND VGND VPWR VPWR registers\[53\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17857_ registers\[16\]\[50\] registers\[17\]\[50\] registers\[18\]\[50\] registers\[19\]\[50\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__mux4_1
XFILLER_26_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_226_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35642_ clknet_leaf_302_CLK _03756_ VGND VGND VPWR VPWR registers\[11\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_16808_ _14613_ VGND VGND VPWR VPWR _15302_ sky130_fd_sc_hd__buf_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32854_ clknet_leaf_65_CLK _00968_ VGND VGND VPWR VPWR registers\[54\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17788_ registers\[28\]\[48\] registers\[29\]\[48\] registers\[30\]\[48\] registers\[31\]\[48\]
+ _04363_ _04364_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux4_1
XFILLER_130_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31805_ registers\[59\]\[59\] net55 _14403_ VGND VGND VPWR VPWR _14413_ sky130_fd_sc_hd__mux2_1
X_19527_ registers\[28\]\[32\] registers\[29\]\[32\] registers\[30\]\[32\] registers\[31\]\[32\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__mux4_1
X_35573_ clknet_leaf_324_CLK _03687_ VGND VGND VPWR VPWR registers\[12\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_16739_ _14991_ _15230_ _15233_ _14996_ VGND VGND VPWR VPWR _15234_ sky130_fd_sc_hd__a22o_1
X_32785_ clknet_leaf_174_CLK _00899_ VGND VGND VPWR VPWR registers\[55\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34524_ clknet_leaf_0_CLK _02638_ VGND VGND VPWR VPWR registers\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19458_ registers\[20\]\[30\] registers\[21\]\[30\] registers\[22\]\[30\] registers\[23\]\[30\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__mux4_1
XFILLER_35_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31736_ registers\[59\]\[26\] net19 _14370_ VGND VGND VPWR VPWR _14377_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18409_ _05122_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__buf_4
XFILLER_195_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34455_ clknet_leaf_87_CLK _02569_ VGND VGND VPWR VPWR registers\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_349_CLK clknet_6_46__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_349_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31667_ _14340_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__clkbuf_1
X_19389_ _05067_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__buf_6
XFILLER_50_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33406_ clknet_leaf_274_CLK _01520_ VGND VGND VPWR VPWR registers\[46\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21420_ registers\[48\]\[21\] registers\[49\]\[21\] registers\[50\]\[21\] registers\[51\]\[21\]
+ _07986_ _07987_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__mux4_1
X_30618_ registers\[12\]\[8\] _12951_ _13780_ VGND VGND VPWR VPWR _13789_ sky130_fd_sc_hd__mux2_1
X_34386_ clknet_leaf_100_CLK _02500_ VGND VGND VPWR VPWR registers\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31598_ _14304_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36125_ clknet_leaf_53_CLK _04239_ VGND VGND VPWR VPWR registers\[49\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33337_ clknet_leaf_280_CLK _01451_ VGND VGND VPWR VPWR registers\[47\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_21351_ registers\[8\]\[19\] registers\[9\]\[19\] registers\[10\]\[19\] registers\[11\]\[19\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__mux4_1
XFILLER_198_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30549_ _13752_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20302_ _07007_ _07010_ _06880_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__o21ba_1
X_24070_ _10211_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36056_ clknet_leaf_52_CLK _04170_ VGND VGND VPWR VPWR registers\[59\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21282_ registers\[12\]\[17\] registers\[13\]\[17\] registers\[14\]\[17\] registers\[15\]\[17\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__mux4_1
X_33268_ clknet_leaf_350_CLK _01382_ VGND VGND VPWR VPWR registers\[48\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35007_ clknet_leaf_306_CLK _03121_ VGND VGND VPWR VPWR registers\[21\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_23021_ _09610_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
X_32219_ clknet_leaf_238_CLK _00333_ VGND VGND VPWR VPWR registers\[9\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_20233_ registers\[28\]\[52\] registers\[29\]\[52\] registers\[30\]\[52\] registers\[31\]\[52\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__mux4_1
XFILLER_116_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33199_ clknet_leaf_378_CLK _01313_ VGND VGND VPWR VPWR registers\[4\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_235_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20164_ registers\[20\]\[50\] registers\[21\]\[50\] registers\[22\]\[50\] registers\[23\]\[50\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__mux4_1
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_226_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27760_ registers\[33\]\[29\] _10365_ _12244_ VGND VGND VPWR VPWR _12254_ sky130_fd_sc_hd__mux2_1
X_20095_ _05051_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__clkbuf_8
X_24972_ _10719_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26711_ registers\[40\]\[11\] _10328_ _11669_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__mux2_1
XFILLER_58_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35909_ clknet_leaf_230_CLK _04023_ VGND VGND VPWR VPWR registers\[7\]\[55\] sky130_fd_sc_hd__dfxtp_1
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ _09598_ registers\[60\]\[40\] _10133_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__mux2_1
X_27691_ _12217_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_217_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_218_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29430_ _09702_ registers\[21\]\[21\] _13162_ VGND VGND VPWR VPWR _13164_ sky130_fd_sc_hd__mux2_1
XFILLER_242_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23854_ _10097_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
X_26642_ _10821_ registers\[41\]\[43\] _11630_ VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__mux2_1
XFILLER_79_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_605 _05102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_616 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _09439_ _09442_ _07369_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__o21ba_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29361_ _13127_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_627 _05122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26573_ _10751_ registers\[41\]\[10\] _11597_ VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__mux2_1
XANTENNA_638 _05152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23785_ _10060_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__clkbuf_1
X_20997_ _07683_ _07686_ _07339_ _07341_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__o211a_1
XANTENNA_649 _05165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28312_ _12544_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_197_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22736_ registers\[52\]\[59\] registers\[53\]\[59\] registers\[54\]\[59\] registers\[55\]\[59\]
+ _07279_ _07282_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__mux4_1
XFILLER_168_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25524_ registers\[4\]\[28\] _10363_ _11034_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__mux2_1
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29292_ _13068_ VGND VGND VPWR VPWR _13091_ sky130_fd_sc_hd__buf_4
XFILLER_129_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28243_ _12508_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__clkbuf_1
X_25455_ _11004_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22667_ _09148_ _09307_ _09308_ _09153_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__a22o_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24406_ _10413_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
X_21618_ _08119_ _08288_ _08289_ _08124_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__a22o_1
X_28174_ _11799_ registers\[30\]\[33\] _12468_ VGND VGND VPWR VPWR _12472_ sky130_fd_sc_hd__mux2_1
X_25386_ _10968_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__clkbuf_1
X_22598_ _09104_ _09241_ _09242_ _09107_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__a22o_1
XFILLER_127_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27125_ _11832_ registers\[38\]\[49\] _11909_ VGND VGND VPWR VPWR _11919_ sky130_fd_sc_hd__mux2_1
X_24337_ _10366_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
X_21549_ registers\[44\]\[25\] registers\[45\]\[25\] registers\[46\]\[25\] registers\[47\]\[25\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__mux4_1
XFILLER_194_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27056_ _11763_ registers\[38\]\[16\] _11876_ VGND VGND VPWR VPWR _11883_ sky130_fd_sc_hd__mux2_1
X_24268_ registers\[57\]\[7\] _10319_ _10305_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__mux2_1
XFILLER_154_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26007_ _10862_ registers\[46\]\[63\] _11229_ VGND VGND VPWR VPWR _11299_ sky130_fd_sc_hd__mux2_1
X_23219_ _09741_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24199_ _09603_ registers\[58\]\[42\] _10277_ VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__mux2_1
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1004 _11832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1015 _12150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1026 _12718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1037 _13139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1048 _13281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18760_ registers\[32\]\[11\] registers\[33\]\[11\] registers\[34\]\[11\] registers\[35\]\[11\]
+ _05437_ _05438_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__mux4_1
X_27958_ registers\[32\]\[59\] _10428_ _12348_ VGND VGND VPWR VPWR _12358_ sky130_fd_sc_hd__mux2_1
XTAP_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1059 _13850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ registers\[24\]\[46\] registers\[25\]\[46\] registers\[26\]\[46\] registers\[27\]\[46\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__mux4_1
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26909_ net21 VGND VGND VPWR VPWR _11788_ sky130_fd_sc_hd__clkbuf_4
XTAP_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ registers\[56\]\[9\] registers\[57\]\[9\] registers\[58\]\[9\] registers\[59\]\[9\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__mux4_1
XFILLER_62_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_5_18_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_18_0_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27889_ registers\[32\]\[26\] _10359_ _12315_ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__mux2_1
XTAP_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17642_ _14564_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__buf_6
XFILLER_212_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29628_ registers\[20\]\[51\] _13042_ _13266_ VGND VGND VPWR VPWR _13268_ sky130_fd_sc_hd__mux2_1
XFILLER_64_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_247_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17573_ _15830_ _04356_ _04357_ _15833_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a22o_1
X_29559_ _13231_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19312_ _05844_ _06047_ _06048_ _05849_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__a22o_1
XFILLER_182_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16524_ _15020_ _15025_ _14959_ VGND VGND VPWR VPWR _15026_ sky130_fd_sc_hd__o21ba_1
XFILLER_189_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32570_ clknet_leaf_304_CLK _00684_ VGND VGND VPWR VPWR registers\[5\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31521_ _09802_ registers\[6\]\[52\] _14261_ VGND VGND VPWR VPWR _14264_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19243_ _05978_ _05981_ _05851_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__o21ba_1
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16455_ _14613_ VGND VGND VPWR VPWR _14959_ sky130_fd_sc_hd__buf_2
XFILLER_182_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_220_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34240_ clknet_leaf_270_CLK _02354_ VGND VGND VPWR VPWR registers\[33\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31452_ _14227_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__clkbuf_1
X_19174_ registers\[28\]\[22\] registers\[29\]\[22\] registers\[30\]\[22\] registers\[31\]\[22\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux4_1
XFILLER_34_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_223_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16386_ _14648_ _14887_ _14890_ _14653_ VGND VGND VPWR VPWR _14891_ sky130_fd_sc_hd__a22o_1
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18125_ registers\[40\]\[59\] registers\[41\]\[59\] registers\[42\]\[59\] registers\[43\]\[59\]
+ _04677_ _04678_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux4_1
XFILLER_129_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30403_ _09762_ registers\[14\]\[34\] _13671_ VGND VGND VPWR VPWR _13676_ sky130_fd_sc_hd__mux2_1
XFILLER_247_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34171_ clknet_leaf_282_CLK _02285_ VGND VGND VPWR VPWR registers\[34\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_31383_ _14191_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33122_ clknet_leaf_45_CLK _01236_ VGND VGND VPWR VPWR registers\[50\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_18056_ registers\[24\]\[56\] registers\[25\]\[56\] registers\[26\]\[56\] registers\[27\]\[56\]
+ _04767_ _04768_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__mux4_1
X_30334_ _09660_ registers\[14\]\[1\] _13638_ VGND VGND VPWR VPWR _13640_ sky130_fd_sc_hd__mux2_1
XANTENNA_1 CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17007_ _14594_ VGND VGND VPWR VPWR _15495_ sky130_fd_sc_hd__buf_4
X_33053_ clknet_leaf_51_CLK _01167_ VGND VGND VPWR VPWR registers\[51\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30265_ registers\[15\]\[33\] _13004_ _13599_ VGND VGND VPWR VPWR _13603_ sky130_fd_sc_hd__mux2_1
XFILLER_67_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32004_ clknet_leaf_28_CLK _00177_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30196_ registers\[15\]\[0\] _12931_ _13566_ VGND VGND VPWR VPWR _13567_ sky130_fd_sc_hd__mux2_1
XFILLER_152_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18958_ registers\[20\]\[16\] registers\[21\]\[16\] registers\[22\]\[16\] registers\[23\]\[16\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__mux4_1
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1560 _11585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1571 _12962_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17909_ registers\[44\]\[52\] registers\[45\]\[52\] registers\[46\]\[52\] registers\[47\]\[52\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__mux4_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1582 _14276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33955_ clknet_leaf_47_CLK _02069_ VGND VGND VPWR VPWR registers\[37\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18889_ _05501_ _05636_ _05637_ _05506_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a22o_1
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1593 _14539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32906_ clknet_leaf_162_CLK _01020_ VGND VGND VPWR VPWR registers\[54\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_20920_ registers\[48\]\[7\] registers\[49\]\[7\] registers\[50\]\[7\] registers\[51\]\[7\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__mux4_1
XFILLER_6_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33886_ clknet_leaf_23_CLK _02000_ VGND VGND VPWR VPWR registers\[38\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_215_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32837_ clknet_leaf_200_CLK _00951_ VGND VGND VPWR VPWR registers\[55\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_20851_ registers\[52\]\[5\] registers\[53\]\[5\] registers\[54\]\[5\] registers\[55\]\[5\]
+ _07332_ _07334_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__mux4_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35625_ clknet_leaf_460_CLK _03739_ VGND VGND VPWR VPWR registers\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23570_ _09946_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35556_ clknet_leaf_467_CLK _03670_ VGND VGND VPWR VPWR registers\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32768_ clknet_leaf_267_CLK _00882_ VGND VGND VPWR VPWR registers\[56\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_20782_ registers\[48\]\[3\] registers\[49\]\[3\] registers\[50\]\[3\] registers\[51\]\[3\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__mux4_1
XFILLER_223_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22521_ registers\[8\]\[52\] registers\[9\]\[52\] registers\[10\]\[52\] registers\[11\]\[52\]
+ _08920_ _08921_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__mux4_1
X_34507_ clknet_leaf_151_CLK _02621_ VGND VGND VPWR VPWR registers\[2\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_31719_ registers\[59\]\[18\] net10 _14359_ VGND VGND VPWR VPWR _14368_ sky130_fd_sc_hd__mux2_1
X_35487_ clknet_leaf_482_CLK _03601_ VGND VGND VPWR VPWR registers\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32699_ clknet_leaf_283_CLK _00813_ VGND VGND VPWR VPWR registers\[57\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_25240_ _10891_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__clkbuf_1
X_34438_ clknet_leaf_213_CLK _02552_ VGND VGND VPWR VPWR registers\[30\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_22452_ _08958_ _09099_ _09100_ _08961_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__a22o_1
XFILLER_210_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21403_ _07315_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__buf_4
X_25171_ net54 VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__clkbuf_8
XFILLER_202_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34369_ clknet_leaf_203_CLK _02483_ VGND VGND VPWR VPWR registers\[31\]\[51\] sky130_fd_sc_hd__dfxtp_1
X_22383_ _08958_ _09030_ _09033_ _08961_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__a22o_1
XFILLER_124_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_36108_ clknet_leaf_167_CLK _04222_ VGND VGND VPWR VPWR registers\[59\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_24122_ _10239_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__clkbuf_1
X_21334_ _08014_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36039_ clknet_leaf_196_CLK _04153_ VGND VGND VPWR VPWR registers\[63\]\[57\] sky130_fd_sc_hd__dfxtp_1
X_28930_ _12869_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__clkbuf_1
X_24053_ _10202_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__clkbuf_1
X_21265_ _07776_ _07945_ _07946_ _07781_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__a22o_1
XFILLER_104_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_50_CLK sky130_fd_sc_hd__clkbuf_16
X_23004_ _09514_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__buf_4
X_20216_ _06776_ _06925_ _06926_ _06782_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__a22o_1
X_28861_ _11811_ registers\[25\]\[39\] _12823_ VGND VGND VPWR VPWR _12833_ sky130_fd_sc_hd__mux2_1
X_21196_ registers\[44\]\[15\] registers\[45\]\[15\] registers\[46\]\[15\] registers\[47\]\[15\]
+ _07706_ _07707_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__mux4_1
XFILLER_46_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27812_ _12281_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__clkbuf_1
X_20147_ _05122_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__buf_4
XFILLER_172_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_217_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28792_ _11742_ registers\[25\]\[6\] _12790_ VGND VGND VPWR VPWR _12797_ sky130_fd_sc_hd__mux2_1
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27743_ _12245_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__clkbuf_1
X_20078_ _06717_ _06791_ _06792_ _06720_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__a22o_1
X_24955_ _10710_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _09582_ registers\[60\]\[32\] _10122_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__mux2_1
X_27674_ registers\[34\]\[52\] _10414_ _12206_ VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__mux2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24886_ _10674_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_402 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29413_ _09685_ registers\[21\]\[13\] _13151_ VGND VGND VPWR VPWR _13155_ sky130_fd_sc_hd__mux2_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26625_ _10804_ registers\[41\]\[35\] _11619_ VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__mux2_1
XFILLER_73_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23837_ _10087_ VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__buf_12
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_424 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_446 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29344_ _13118_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_457 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26556_ _10735_ registers\[41\]\[2\] _11586_ VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__mux2_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23768_ _09580_ registers\[29\]\[31\] _10050_ VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__mux2_1
XANTENNA_468 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_479 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_207_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25507_ _11011_ VGND VGND VPWR VPWR _11034_ sky130_fd_sc_hd__buf_4
X_22719_ registers\[28\]\[58\] registers\[29\]\[58\] registers\[30\]\[58\] registers\[31\]\[58\]
+ _09178_ _09179_ VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__mux4_1
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29275_ _13082_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__clkbuf_1
X_23699_ _09651_ _10013_ VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__nor2_8
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26487_ _10802_ registers\[42\]\[34\] _11547_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__mux2_1
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16240_ registers\[40\]\[5\] registers\[41\]\[5\] registers\[42\]\[5\] registers\[43\]\[5\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14749_ sky130_fd_sc_hd__mux4_1
X_28226_ _11851_ registers\[30\]\[58\] _12490_ VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__mux2_1
XFILLER_185_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25438_ _10842_ registers\[50\]\[53\] _10992_ VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__mux2_1
XFILLER_185_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_1336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16171_ _14677_ _14682_ _14614_ VGND VGND VPWR VPWR _14683_ sky130_fd_sc_hd__o21ba_1
XFILLER_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28157_ _11782_ registers\[30\]\[25\] _12457_ VGND VGND VPWR VPWR _12463_ sky130_fd_sc_hd__mux2_1
X_25369_ _10772_ registers\[50\]\[20\] _10959_ VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__mux2_1
XFILLER_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27108_ _11910_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28088_ _12426_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19930_ registers\[60\]\[44\] registers\[61\]\[44\] registers\[62\]\[44\] registers\[63\]\[44\]
+ _06648_ _06442_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__mux4_1
XFILLER_99_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27039_ _11746_ registers\[38\]\[8\] _11865_ VGND VGND VPWR VPWR _11874_ sky130_fd_sc_hd__mux2_1
XFILLER_181_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_41_CLK sky130_fd_sc_hd__clkbuf_16
X_30050_ _13489_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19861_ registers\[56\]\[42\] registers\[57\]\[42\] registers\[58\]\[42\] registers\[59\]\[42\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__mux4_1
XFILLER_134_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_5_1_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_1_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_110_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18812_ registers\[12\]\[12\] registers\[13\]\[12\] registers\[14\]\[12\] registers\[15\]\[12\]
+ _05251_ _05252_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__mux4_1
XTAP_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput93 net93 VGND VGND VPWR VPWR D1[12] sky130_fd_sc_hd__buf_2
XFILLER_231_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19792_ registers\[8\]\[40\] registers\[9\]\[40\] registers\[10\]\[40\] registers\[11\]\[40\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__mux4_1
XFILLER_228_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18743_ _05136_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__clkbuf_4
XTAP_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33740_ clknet_leaf_171_CLK _01854_ VGND VGND VPWR VPWR registers\[41\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_18674_ registers\[16\]\[8\] registers\[17\]\[8\] registers\[18\]\[8\] registers\[19\]\[8\]
+ _05357_ _05358_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__mux4_1
XFILLER_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30952_ _13964_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__clkbuf_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _14529_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__buf_6
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33671_ clknet_leaf_243_CLK _01785_ VGND VGND VPWR VPWR registers\[42\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_184_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30883_ _13928_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35410_ clknet_leaf_77_CLK _03524_ VGND VGND VPWR VPWR registers\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32622_ clknet_leaf_371_CLK _00736_ VGND VGND VPWR VPWR registers\[58\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_17556_ registers\[44\]\[42\] registers\[45\]\[42\] registers\[46\]\[42\] registers\[47\]\[42\]
+ _15950_ _15951_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__mux4_1
XANTENNA_980 _11229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35341_ clknet_leaf_148_CLK _03455_ VGND VGND VPWR VPWR registers\[16\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16507_ _14863_ _15007_ _15008_ _14867_ VGND VGND VPWR VPWR _15009_ sky130_fd_sc_hd__a22o_1
XFILLER_60_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_991 _11729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32553_ clknet_leaf_401_CLK _00667_ VGND VGND VPWR VPWR registers\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17487_ registers\[52\]\[40\] registers\[53\]\[40\] registers\[54\]\[40\] registers\[55\]\[40\]
+ _15820_ _15821_ VGND VGND VPWR VPWR _15961_ sky130_fd_sc_hd__mux4_1
X_31504_ _09784_ registers\[6\]\[44\] _14250_ VGND VGND VPWR VPWR _14255_ sky130_fd_sc_hd__mux2_1
XFILLER_20_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19226_ _05755_ _05963_ _05964_ _05759_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a22o_1
X_35272_ clknet_leaf_153_CLK _03386_ VGND VGND VPWR VPWR registers\[17\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_16438_ registers\[12\]\[10\] registers\[13\]\[10\] registers\[14\]\[10\] registers\[15\]\[10\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14942_ sky130_fd_sc_hd__mux4_1
X_32484_ clknet_leaf_446_CLK _00598_ VGND VGND VPWR VPWR registers\[60\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_34223_ clknet_leaf_355_CLK _02337_ VGND VGND VPWR VPWR registers\[33\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31435_ _09681_ registers\[6\]\[11\] _14217_ VGND VGND VPWR VPWR _14219_ sky130_fd_sc_hd__mux2_1
X_19157_ _05747_ _05896_ _05897_ _05753_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__a22o_1
X_16369_ _14578_ VGND VGND VPWR VPWR _14875_ sky130_fd_sc_hd__buf_4
XFILLER_157_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ _04873_ _04876_ _04619_ _04620_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__o211a_1
X_34154_ clknet_leaf_431_CLK _02268_ VGND VGND VPWR VPWR registers\[34\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31366_ _14182_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__clkbuf_1
X_19088_ _05113_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_121_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33105_ clknet_leaf_74_CLK _01219_ VGND VGND VPWR VPWR registers\[50\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30317_ registers\[15\]\[58\] _13056_ _13621_ VGND VGND VPWR VPWR _13630_ sky130_fd_sc_hd__mux2_1
X_18039_ registers\[36\]\[56\] registers\[37\]\[56\] registers\[38\]\[56\] registers\[39\]\[56\]
+ _04506_ _04507_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__mux4_1
XFILLER_195_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34085_ clknet_leaf_433_CLK _02199_ VGND VGND VPWR VPWR registers\[35\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_31297_ _14134_ VGND VGND VPWR VPWR _14146_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_32_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_32_CLK sky130_fd_sc_hd__clkbuf_16
X_33036_ clknet_leaf_142_CLK _01150_ VGND VGND VPWR VPWR registers\[52\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21050_ _07315_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__buf_4
XFILLER_67_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30248_ registers\[15\]\[25\] _12987_ _13588_ VGND VGND VPWR VPWR _13594_ sky130_fd_sc_hd__mux2_1
XFILLER_154_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20001_ registers\[8\]\[46\] registers\[9\]\[46\] registers\[10\]\[46\] registers\[11\]\[46\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__mux4_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30179_ _13557_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1390 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34987_ clknet_leaf_458_CLK _03101_ VGND VGND VPWR VPWR registers\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24740_ _10597_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
X_21952_ _07295_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__buf_4
X_33938_ clknet_leaf_120_CLK _02052_ VGND VGND VPWR VPWR registers\[37\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20903_ _07373_ _07592_ _07595_ _07383_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__a22o_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24671_ _10560_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
X_33869_ clknet_leaf_147_CLK _01983_ VGND VGND VPWR VPWR registers\[3\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_21883_ _08267_ _08546_ _08547_ _08270_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_99_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_99_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26410_ _10860_ registers\[43\]\[62\] _11442_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__mux2_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23622_ _09973_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
X_20834_ registers\[28\]\[4\] registers\[29\]\[4\] registers\[30\]\[4\] registers\[31\]\[4\]
+ _07463_ _07464_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__mux4_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35608_ clknet_leaf_15_CLK _03722_ VGND VGND VPWR VPWR registers\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_27390_ _12058_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_223_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23553_ _09640_ registers\[19\]\[60\] _09869_ VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__mux2_1
XFILLER_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26341_ _10791_ registers\[43\]\[29\] _11465_ VGND VGND VPWR VPWR _11475_ sky130_fd_sc_hd__mux2_1
X_20765_ _07373_ _07460_ _07461_ _07383_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__a22o_1
X_35539_ clknet_leaf_79_CLK _03653_ VGND VGND VPWR VPWR registers\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22504_ registers\[40\]\[52\] registers\[41\]\[52\] registers\[42\]\[52\] registers\[43\]\[52\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__mux4_1
XFILLER_211_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26272_ _11438_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
X_29060_ _12940_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1047 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23484_ _09571_ registers\[19\]\[27\] _09892_ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1000 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20696_ _07300_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__buf_12
XFILLER_149_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25223_ _10882_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__clkbuf_1
X_28011_ _12363_ VGND VGND VPWR VPWR _12386_ sky130_fd_sc_hd__buf_4
X_22435_ _09077_ _09082_ _09083_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__o21ba_1
XFILLER_241_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25154_ _10840_ registers\[52\]\[52\] _10836_ VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__mux2_1
X_22366_ registers\[48\]\[48\] registers\[49\]\[48\] registers\[50\]\[48\] registers\[51\]\[48\]
+ _09015_ _09016_ VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__mux4_1
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24105_ _10229_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21317_ registers\[8\]\[18\] registers\[9\]\[18\] registers\[10\]\[18\] registers\[11\]\[18\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__mux4_1
XFILLER_151_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29962_ _13443_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__clkbuf_1
X_25085_ _10730_ VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__clkbuf_8
X_22297_ registers\[52\]\[46\] registers\[53\]\[46\] registers\[54\]\[46\] registers\[55\]\[46\]
+ _08948_ _08949_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__mux4_1
XFILLER_184_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_23_CLK sky130_fd_sc_hd__clkbuf_16
X_28913_ _09651_ _10013_ _11084_ VGND VGND VPWR VPWR _12860_ sky130_fd_sc_hd__nor3_4
XFILLER_190_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24036_ _10193_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21248_ registers\[4\]\[16\] registers\[5\]\[16\] registers\[6\]\[16\] registers\[7\]\[16\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__mux4_1
XFILLER_105_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29893_ registers\[18\]\[49\] _13037_ _13397_ VGND VGND VPWR VPWR _13407_ sky130_fd_sc_hd__mux2_1
XFILLER_77_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28844_ _12824_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__clkbuf_1
X_21179_ registers\[4\]\[14\] registers\[5\]\[14\] registers\[6\]\[14\] registers\[7\]\[14\]
+ _07659_ _07660_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__mux4_1
XFILLER_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28775_ _12787_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25987_ _10842_ registers\[46\]\[53\] _11285_ VGND VGND VPWR VPWR _11289_ sky130_fd_sc_hd__mux2_1
XFILLER_24_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27726_ _12236_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__clkbuf_1
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24938_ _10701_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27657_ registers\[34\]\[44\] _10397_ _12195_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__mux2_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24869_ _10665_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__clkbuf_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_221 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17410_ registers\[56\]\[38\] registers\[57\]\[38\] registers\[58\]\[38\] registers\[59\]\[38\]
+ _15752_ _15885_ VGND VGND VPWR VPWR _15886_ sky130_fd_sc_hd__mux4_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26608_ _10787_ registers\[41\]\[27\] _11608_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__mux2_1
XFILLER_57_1220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__buf_4
XANTENNA_254 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27588_ registers\[34\]\[11\] _10328_ _12162_ VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__mux2_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_276 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29327_ _13109_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__clkbuf_1
X_17341_ registers\[60\]\[36\] registers\[61\]\[36\] registers\[62\]\[36\] registers\[63\]\[36\]
+ _15756_ _15550_ VGND VGND VPWR VPWR _15819_ sky130_fd_sc_hd__mux4_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26539_ _10854_ registers\[42\]\[59\] _11569_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__mux2_1
XFILLER_186_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_298 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_1166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29258_ _13073_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__clkbuf_1
X_17272_ _14529_ VGND VGND VPWR VPWR _15752_ sky130_fd_sc_hd__buf_6
XFILLER_140_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19011_ _05092_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__clkbuf_4
X_28209_ _12434_ VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__buf_4
XFILLER_174_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16223_ registers\[0\]\[4\] registers\[1\]\[4\] registers\[2\]\[4\] registers\[3\]\[4\]
+ _14563_ _14565_ VGND VGND VPWR VPWR _14733_ sky130_fd_sc_hd__mux4_1
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29189_ registers\[23\]\[44\] _13027_ _13019_ VGND VGND VPWR VPWR _13028_ sky130_fd_sc_hd__mux2_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31220_ _14105_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__clkbuf_1
X_16154_ _14540_ _14664_ _14665_ _14551_ VGND VGND VPWR VPWR _14666_ sky130_fd_sc_hd__a22o_1
XFILLER_127_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31151_ _14069_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16085_ _14588_ _14591_ _14596_ _14598_ VGND VGND VPWR VPWR _14599_ sky130_fd_sc_hd__a22o_1
XFILLER_177_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_14_CLK sky130_fd_sc_hd__clkbuf_16
X_30102_ _13494_ VGND VGND VPWR VPWR _13517_ sky130_fd_sc_hd__buf_4
XFILLER_68_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1040 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19913_ registers\[20\]\[43\] registers\[21\]\[43\] registers\[22\]\[43\] registers\[23\]\[43\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__mux4_1
X_31082_ registers\[0\]\[36\] _13010_ _14026_ VGND VGND VPWR VPWR _14033_ sky130_fd_sc_hd__mux2_1
XFILLER_190_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30033_ registers\[17\]\[51\] _13042_ _13479_ VGND VGND VPWR VPWR _13481_ sky130_fd_sc_hd__mux2_1
XFILLER_151_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19844_ _06530_ _06564_ _06565_ _06535_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__a22o_1
X_34910_ clknet_leaf_491_CLK _03024_ VGND VGND VPWR VPWR registers\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35890_ clknet_leaf_379_CLK _04004_ VGND VGND VPWR VPWR registers\[7\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34841_ clknet_leaf_4_CLK _02955_ VGND VGND VPWR VPWR registers\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_19775_ _06226_ _06496_ _06497_ _06231_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__a22o_1
X_16987_ _15198_ _15473_ _15474_ _15204_ VGND VGND VPWR VPWR _15475_ sky130_fd_sc_hd__a22o_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18726_ _05404_ _05477_ _05478_ _05410_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__a22o_1
XFILLER_83_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34772_ clknet_leaf_88_CLK _02886_ VGND VGND VPWR VPWR registers\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31984_ clknet_leaf_21_CLK _00155_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33723_ clknet_leaf_279_CLK _01837_ VGND VGND VPWR VPWR registers\[41\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_18657_ _05088_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__buf_4
X_30935_ registers\[10\]\[30\] _12997_ _13955_ VGND VGND VPWR VPWR _13956_ sky130_fd_sc_hd__mux2_1
XFILLER_18_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17608_ _04386_ _04391_ _15974_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__o21ba_1
XFILLER_18_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_992 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33654_ clknet_leaf_341_CLK _01768_ VGND VGND VPWR VPWR registers\[42\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1099 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30866_ _09823_ registers\[11\]\[62\] _13850_ VGND VGND VPWR VPWR _13919_ sky130_fd_sc_hd__mux2_1
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18588_ _05039_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__buf_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32605_ clknet_leaf_51_CLK _00719_ VGND VGND VPWR VPWR registers\[58\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ registers\[24\]\[41\] registers\[25\]\[41\] registers\[26\]\[41\] registers\[27\]\[41\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__mux4_1
XFILLER_36_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33585_ clknet_leaf_347_CLK _01699_ VGND VGND VPWR VPWR registers\[43\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_189_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30797_ _09751_ registers\[11\]\[29\] _13873_ VGND VGND VPWR VPWR _13883_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35324_ clknet_leaf_189_CLK _03438_ VGND VGND VPWR VPWR registers\[16\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_20550_ _05089_ _07248_ _07249_ _05100_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__a22o_1
X_32536_ clknet_leaf_474_CLK _00650_ VGND VGND VPWR VPWR registers\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19209_ _05945_ _05948_ _05851_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__o21ba_1
X_35255_ clknet_leaf_311_CLK _03369_ VGND VGND VPWR VPWR registers\[17\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_20481_ _05119_ _07182_ _07183_ _05131_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__a22o_1
X_32467_ clknet_leaf_182_CLK _00581_ VGND VGND VPWR VPWR registers\[60\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22220_ _08805_ _08873_ _08874_ _08810_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__a22o_1
XFILLER_121_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34206_ clknet_leaf_22_CLK _02320_ VGND VGND VPWR VPWR registers\[33\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_31418_ _09664_ registers\[6\]\[3\] _14206_ VGND VGND VPWR VPWR _14210_ sky130_fd_sc_hd__mux2_1
X_35186_ clknet_leaf_417_CLK _03300_ VGND VGND VPWR VPWR registers\[18\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32398_ clknet_leaf_109_CLK _00512_ VGND VGND VPWR VPWR registers\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_34137_ clknet_leaf_91_CLK _02251_ VGND VGND VPWR VPWR registers\[34\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_22151_ registers\[40\]\[42\] registers\[41\]\[42\] registers\[42\]\[42\] registers\[43\]\[42\]
+ _08806_ _08807_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__mux4_1
XFILLER_121_1097 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31349_ _14173_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21102_ registers\[56\]\[12\] registers\[57\]\[12\] registers\[58\]\[12\] registers\[59\]\[12\]
+ _07508_ _07641_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__mux4_1
XTAP_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34068_ clknet_leaf_121_CLK _02182_ VGND VGND VPWR VPWR registers\[35\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22082_ _08734_ _08739_ _08740_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__o21ba_1
XTAP_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_1173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33019_ clknet_leaf_286_CLK _01133_ VGND VGND VPWR VPWR registers\[52\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_21033_ registers\[8\]\[10\] registers\[9\]\[10\] registers\[10\]\[10\] registers\[11\]\[10\]
+ _07548_ _07549_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__mux4_1
XFILLER_99_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25910_ _11248_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_232_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26890_ _11775_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25841_ _10831_ registers\[47\]\[48\] _11203_ VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_214_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28560_ _11780_ registers\[27\]\[24\] _12670_ VGND VGND VPWR VPWR _12675_ sky130_fd_sc_hd__mux2_1
X_25772_ _10762_ registers\[47\]\[15\] _11170_ VGND VGND VPWR VPWR _11176_ sky130_fd_sc_hd__mux2_1
X_22984_ _09585_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_216_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27511_ _12077_ VGND VGND VPWR VPWR _12122_ sky130_fd_sc_hd__buf_4
X_24723_ _09517_ registers\[54\]\[1\] _10587_ VGND VGND VPWR VPWR _10589_ sky130_fd_sc_hd__mux2_1
X_28491_ _12638_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21935_ registers\[36\]\[36\] registers\[37\]\[36\] registers\[38\]\[36\] registers\[39\]\[36\]
+ _08292_ _08293_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__mux4_1
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27442_ _11744_ registers\[35\]\[7\] _12078_ VGND VGND VPWR VPWR _12086_ sky130_fd_sc_hd__mux2_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24654_ _10551_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
X_21866_ registers\[32\]\[34\] registers\[33\]\[34\] registers\[34\]\[34\] registers\[35\]\[34\]
+ _08359_ _08360_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__mux4_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _07326_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__buf_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _09964_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
X_27373_ _12049_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24585_ _10515_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21797_ _07281_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29112_ _12975_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26324_ _11466_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__clkbuf_1
X_23536_ _09927_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
X_20748_ _07439_ _07444_ _07310_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__o21ba_1
XFILLER_141_1418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29043_ _12928_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26255_ _10840_ registers\[44\]\[52\] _11427_ VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__mux2_1
XFILLER_195_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23467_ _09554_ registers\[19\]\[19\] _09881_ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__mux2_1
XFILLER_52_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20679_ _07377_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__buf_6
XFILLER_52_1172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22418_ registers\[16\]\[49\] registers\[17\]\[49\] registers\[18\]\[49\] registers\[19\]\[49\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__mux4_1
X_25206_ _10873_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23398_ _09853_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
X_26186_ _11393_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25137_ net42 VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__buf_2
X_22349_ registers\[20\]\[47\] registers\[21\]\[47\] registers\[22\]\[47\] registers\[23\]\[47\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__mux4_1
XFILLER_178_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29945_ _13434_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25068_ _10782_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24019_ _09559_ registers\[5\]\[21\] _10183_ VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__mux2_1
X_16910_ _15377_ _15384_ _15393_ _15400_ VGND VGND VPWR VPWR _15401_ sky130_fd_sc_hd__or4_4
XFILLER_105_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17890_ _04486_ _04664_ _04665_ _04489_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__a22o_1
X_29876_ _13398_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28827_ _12815_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__clkbuf_1
X_16841_ _15333_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19560_ registers\[20\]\[33\] registers\[21\]\[33\] registers\[22\]\[33\] registers\[23\]\[33\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux4_1
XFILLER_8_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28758_ _11843_ registers\[26\]\[54\] _12774_ VGND VGND VPWR VPWR _12779_ sky130_fd_sc_hd__mux2_1
X_16772_ registers\[44\]\[20\] registers\[45\]\[20\] registers\[46\]\[20\] registers\[47\]\[20\]
+ _15264_ _15265_ VGND VGND VPWR VPWR _15266_ sky130_fd_sc_hd__mux4_2
XFILLER_115_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_247_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_225_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_219_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18511_ _05204_ _05268_ _05269_ _05207_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__a22o_1
XFILLER_92_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_1022 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27709_ _12227_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19491_ _06187_ _06221_ _06222_ _06192_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__a22o_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28689_ _11774_ registers\[26\]\[21\] _12741_ VGND VGND VPWR VPWR _12743_ sky130_fd_sc_hd__mux2_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _05197_ _05200_ _05201_ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__a22o_1
X_30720_ _13842_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__clkbuf_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_CLK clknet_6_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_3_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _05038_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__buf_12
X_30651_ _13806_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__clkbuf_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17324_ _15633_ _15801_ _15802_ _15636_ VGND VGND VPWR VPWR _15803_ sky130_fd_sc_hd__a22o_1
XFILLER_144_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33370_ clknet_leaf_32_CLK _01484_ VGND VGND VPWR VPWR registers\[46\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_30582_ _09808_ registers\[13\]\[55\] _13764_ VGND VGND VPWR VPWR _13770_ sky130_fd_sc_hd__mux2_1
XFILLER_187_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1026 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32321_ clknet_leaf_221_CLK _00435_ VGND VGND VPWR VPWR registers\[19\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17255_ _15730_ _15735_ _15631_ VGND VGND VPWR VPWR _15736_ sky130_fd_sc_hd__o21ba_1
XFILLER_70_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16206_ registers\[40\]\[4\] registers\[41\]\[4\] registers\[42\]\[4\] registers\[43\]\[4\]
+ _14649_ _14650_ VGND VGND VPWR VPWR _14716_ sky130_fd_sc_hd__mux4_1
X_35040_ clknet_leaf_489_CLK _03154_ VGND VGND VPWR VPWR registers\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_32252_ clknet_leaf_282_CLK _00366_ VGND VGND VPWR VPWR registers\[39\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17186_ registers\[24\]\[31\] registers\[25\]\[31\] registers\[26\]\[31\] registers\[27\]\[31\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15669_ sky130_fd_sc_hd__mux4_1
Xclkbuf_6_50__f_CLK clknet_5_25_0_CLK VGND VGND VPWR VPWR clknet_6_50__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31203_ _14096_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__clkbuf_1
X_16137_ _14493_ VGND VGND VPWR VPWR _14649_ sky130_fd_sc_hd__buf_6
XFILLER_31_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32183_ clknet_leaf_486_CLK _00297_ VGND VGND VPWR VPWR registers\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31134_ registers\[0\]\[61\] _13062_ _13992_ VGND VGND VPWR VPWR _14060_ sky130_fd_sc_hd__mux2_1
XFILLER_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16068_ _14581_ VGND VGND VPWR VPWR _14582_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35942_ clknet_leaf_456_CLK _04056_ VGND VGND VPWR VPWR registers\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_31065_ registers\[0\]\[28\] _12993_ _14015_ VGND VGND VPWR VPWR _14024_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1076 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30016_ registers\[17\]\[43\] _13025_ _13468_ VGND VGND VPWR VPWR _13472_ sky130_fd_sc_hd__mux2_1
XFILLER_110_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19827_ _06433_ _06547_ _06548_ _06439_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__a22o_1
X_35873_ clknet_leaf_481_CLK _03987_ VGND VGND VPWR VPWR registers\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_34824_ clknet_leaf_219_CLK _02938_ VGND VGND VPWR VPWR registers\[24\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_19758_ registers\[0\]\[39\] registers\[1\]\[39\] registers\[2\]\[39\] registers\[3\]\[39\]
+ _06173_ _06174_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__mux4_1
XFILLER_204_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_237_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18709_ registers\[20\]\[9\] registers\[21\]\[9\] registers\[22\]\[9\] registers\[23\]\[9\]
+ _05155_ _05157_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__mux4_1
X_34755_ clknet_leaf_224_CLK _02869_ VGND VGND VPWR VPWR registers\[25\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19689_ registers\[4\]\[37\] registers\[5\]\[37\] registers\[6\]\[37\] registers\[7\]\[37\]
+ _06109_ _06110_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__mux4_1
X_31967_ clknet_leaf_4_CLK _00136_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
XFILLER_224_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21720_ registers\[40\]\[30\] registers\[41\]\[30\] registers\[42\]\[30\] registers\[43\]\[30\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__mux4_1
XFILLER_227_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30918_ registers\[10\]\[22\] _12981_ _13944_ VGND VGND VPWR VPWR _13947_ sky130_fd_sc_hd__mux2_1
X_33706_ clknet_leaf_428_CLK _01820_ VGND VGND VPWR VPWR registers\[41\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_224_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34686_ clknet_leaf_179_CLK _02800_ VGND VGND VPWR VPWR registers\[26\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31898_ _09773_ registers\[49\]\[39\] _14452_ VGND VGND VPWR VPWR _14462_ sky130_fd_sc_hd__mux2_1
XFILLER_212_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21651_ registers\[44\]\[28\] registers\[45\]\[28\] registers\[46\]\[28\] registers\[47\]\[28\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__mux4_1
XFILLER_75_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33637_ clknet_leaf_57_CLK _01751_ VGND VGND VPWR VPWR registers\[42\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_30849_ _13910_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_887 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_244_1453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_220_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20602_ _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__buf_12
XFILLER_21_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24370_ _10304_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__buf_4
XFILLER_127_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21582_ registers\[36\]\[26\] registers\[37\]\[26\] registers\[38\]\[26\] registers\[39\]\[26\]
+ _07949_ _07950_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__mux4_1
X_33568_ clknet_leaf_32_CLK _01682_ VGND VGND VPWR VPWR registers\[43\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23321_ _09809_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
X_20533_ registers\[4\]\[62\] registers\[5\]\[62\] registers\[6\]\[62\] registers\[7\]\[62\]
+ _05138_ _05139_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__mux4_1
X_32519_ clknet_leaf_198_CLK _00633_ VGND VGND VPWR VPWR registers\[60\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35307_ clknet_leaf_410_CLK _03421_ VGND VGND VPWR VPWR registers\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_948 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33499_ clknet_leaf_31_CLK _01613_ VGND VGND VPWR VPWR registers\[44\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26040_ _10760_ registers\[45\]\[14\] _11312_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__mux2_1
X_23252_ _09763_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
X_20464_ _05136_ _07165_ _07166_ _05146_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a22o_1
X_35238_ clknet_leaf_449_CLK _03352_ VGND VGND VPWR VPWR registers\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22203_ _07303_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__buf_6
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23183_ _09721_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
X_35169_ clknet_leaf_2_CLK _03283_ VGND VGND VPWR VPWR registers\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_20395_ registers\[40\]\[58\] registers\[41\]\[58\] registers\[42\]\[58\] registers\[43\]\[58\]
+ _06913_ _06914_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__mux4_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22134_ _08610_ _08790_ _08791_ _08613_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__a22o_1
XFILLER_134_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27991_ _11750_ registers\[31\]\[10\] _12375_ VGND VGND VPWR VPWR _12376_ sky130_fd_sc_hd__mux2_1
XTAP_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput250 net250 VGND VGND VPWR VPWR D3[39] sky130_fd_sc_hd__buf_2
Xoutput261 net261 VGND VGND VPWR VPWR D3[49] sky130_fd_sc_hd__buf_2
XFILLER_47_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput272 net272 VGND VGND VPWR VPWR D3[59] sky130_fd_sc_hd__buf_2
X_29730_ _13321_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__clkbuf_1
XTAP_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26942_ _11810_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_1
X_22065_ registers\[16\]\[39\] registers\[17\]\[39\] registers\[18\]\[39\] registers\[19\]\[39\]
+ _08622_ _08623_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__mux4_1
XTAP_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21016_ _07433_ _07703_ _07704_ _07438_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__a22o_1
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29661_ _13285_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__clkbuf_1
XTAP_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26873_ _11763_ registers\[3\]\[16\] _11751_ VGND VGND VPWR VPWR _11764_ sky130_fd_sc_hd__mux2_1
XFILLER_248_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28612_ _11832_ registers\[27\]\[49\] _12692_ VGND VGND VPWR VPWR _12702_ sky130_fd_sc_hd__mux2_1
XFILLER_134_1288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25824_ _11158_ VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__buf_4
XFILLER_229_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29592_ registers\[20\]\[34\] _13006_ _13244_ VGND VGND VPWR VPWR _13249_ sky130_fd_sc_hd__mux2_1
XFILLER_207_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28543_ _11763_ registers\[27\]\[16\] _12659_ VGND VGND VPWR VPWR _12666_ sky130_fd_sc_hd__mux2_1
X_25755_ _10745_ registers\[47\]\[7\] _11159_ VGND VGND VPWR VPWR _11167_ sky130_fd_sc_hd__mux2_1
XFILLER_210_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22967_ _09573_ registers\[62\]\[28\] _09557_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__mux2_1
XFILLER_74_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24706_ _10578_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28474_ _12629_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__clkbuf_1
X_21918_ registers\[12\]\[35\] registers\[13\]\[35\] registers\[14\]\[35\] registers\[15\]\[35\]
+ _08516_ _08517_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__mux4_1
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25686_ _11129_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
X_22898_ net61 VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_230_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27425_ _12076_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24637_ _10542_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__clkbuf_1
X_21849_ _08267_ _08513_ _08514_ _08270_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__a22o_1
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_212_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27356_ registers\[36\]\[30\] _10367_ _12040_ VGND VGND VPWR VPWR _12041_ sky130_fd_sc_hd__mux2_1
XFILLER_196_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24568_ _10504_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26307_ _11457_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
X_23519_ _09918_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__clkbuf_1
X_27287_ _11859_ registers\[37\]\[62\] _11935_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24499_ _10468_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
X_29026_ registers\[24\]\[53\] _10416_ _12916_ VGND VGND VPWR VPWR _12920_ sky130_fd_sc_hd__mux2_1
X_17040_ registers\[16\]\[27\] registers\[17\]\[27\] registers\[18\]\[27\] registers\[19\]\[27\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15527_ sky130_fd_sc_hd__mux4_1
XFILLER_99_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26238_ _10823_ registers\[44\]\[44\] _11416_ VGND VGND VPWR VPWR _11421_ sky130_fd_sc_hd__mux2_1
XFILLER_221_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26169_ _10754_ registers\[44\]\[11\] _11383_ VGND VGND VPWR VPWR _11385_ sky130_fd_sc_hd__mux2_1
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18991_ _05501_ _05735_ _05736_ _05506_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a22o_1
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ registers\[44\]\[53\] registers\[45\]\[53\] registers\[46\]\[53\] registers\[47\]\[53\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__mux4_1
XFILLER_124_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29928_ registers\[17\]\[1\] _12937_ _13424_ VGND VGND VPWR VPWR _13426_ sky130_fd_sc_hd__mux2_1
XFILLER_140_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17873_ _04333_ _04647_ _04648_ _04338_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__a22o_1
XFILLER_152_1355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29859_ _13389_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19612_ _06336_ _06339_ _06169_ _06170_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__o211a_1
X_16824_ _15206_ _15315_ _15316_ _15210_ VGND VGND VPWR VPWR _15317_ sky130_fd_sc_hd__a22o_1
X_32870_ clknet_leaf_438_CLK _00984_ VGND VGND VPWR VPWR registers\[54\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31821_ _09662_ registers\[49\]\[2\] _14419_ VGND VGND VPWR VPWR _14422_ sky130_fd_sc_hd__mux2_1
X_19543_ registers\[60\]\[33\] registers\[61\]\[33\] registers\[62\]\[33\] registers\[63\]\[33\]
+ _05962_ _06099_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__mux4_1
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16755_ registers\[4\]\[19\] registers\[5\]\[19\] registers\[6\]\[19\] registers\[7\]\[19\]
+ _15217_ _15218_ VGND VGND VPWR VPWR _15250_ sky130_fd_sc_hd__mux4_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34540_ clknet_leaf_402_CLK _02654_ VGND VGND VPWR VPWR registers\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_19474_ _06090_ _06204_ _06205_ _06096_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__a22o_1
X_31752_ _14385_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16686_ registers\[24\]\[17\] registers\[25\]\[17\] registers\[26\]\[17\] registers\[27\]\[17\]
+ _15082_ _15083_ VGND VGND VPWR VPWR _15183_ sky130_fd_sc_hd__mux4_1
X_18425_ _05119_ _05185_ _05186_ _05131_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a22o_1
XFILLER_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30703_ _13833_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34471_ clknet_leaf_459_CLK _02585_ VGND VGND VPWR VPWR registers\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31683_ _14349_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33422_ clknet_leaf_147_CLK _01536_ VGND VGND VPWR VPWR registers\[45\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_36210_ clknet_leaf_115_CLK _00093_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dfxtp_1
X_18356_ _05059_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30634_ _13797_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17307_ registers\[48\]\[35\] registers\[49\]\[35\] registers\[50\]\[35\] registers\[51\]\[35\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15786_ sky130_fd_sc_hd__mux4_1
X_36141_ clknet_leaf_379_CLK _04255_ VGND VGND VPWR VPWR registers\[49\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_33353_ clknet_leaf_254_CLK _01467_ VGND VGND VPWR VPWR registers\[47\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18287_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30565_ _09791_ registers\[13\]\[47\] _13753_ VGND VGND VPWR VPWR _13761_ sky130_fd_sc_hd__mux2_1
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32304_ clknet_leaf_393_CLK _00418_ VGND VGND VPWR VPWR registers\[19\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_17238_ _15684_ _15717_ _15718_ _15687_ VGND VGND VPWR VPWR _15719_ sky130_fd_sc_hd__a22o_1
X_36072_ clknet_leaf_436_CLK _04186_ VGND VGND VPWR VPWR registers\[59\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_33284_ clknet_leaf_260_CLK _01398_ VGND VGND VPWR VPWR registers\[48\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30496_ _09687_ registers\[13\]\[14\] _13720_ VGND VGND VPWR VPWR _13725_ sky130_fd_sc_hd__mux2_1
X_35023_ clknet_leaf_116_CLK _03137_ VGND VGND VPWR VPWR registers\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32235_ clknet_leaf_424_CLK _00349_ VGND VGND VPWR VPWR registers\[39\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_17169_ registers\[36\]\[31\] registers\[37\]\[31\] registers\[38\]\[31\] registers\[39\]\[31\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15652_ sky130_fd_sc_hd__mux4_1
XFILLER_200_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32166_ clknet_leaf_136_CLK _00280_ VGND VGND VPWR VPWR registers\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_20180_ _06776_ _06890_ _06891_ _06782_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__a22o_1
XFILLER_157_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31117_ _14051_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_233_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32097_ clknet_leaf_484_CLK _00010_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dfxtp_1
XFILLER_97_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35925_ clknet_leaf_78_CLK _04039_ VGND VGND VPWR VPWR registers\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_31048_ _13992_ VGND VGND VPWR VPWR _14015_ sky130_fd_sc_hd__buf_4
XFILLER_233_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35856_ clknet_leaf_107_CLK _03970_ VGND VGND VPWR VPWR registers\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23870_ _09546_ registers\[60\]\[15\] _10100_ VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__mux2_1
XFILLER_226_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22821_ _09454_ _09457_ _07309_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__o21ba_1
X_34807_ clknet_leaf_314_CLK _02921_ VGND VGND VPWR VPWR registers\[24\]\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35787_ clknet_leaf_151_CLK _03901_ VGND VGND VPWR VPWR registers\[0\]\[61\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_809 _09043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32999_ clknet_leaf_437_CLK _01113_ VGND VGND VPWR VPWR registers\[52\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25540_ _11051_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__clkbuf_1
X_22752_ _09388_ _09391_ _09116_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__o21ba_1
X_34738_ clknet_leaf_412_CLK _02852_ VGND VGND VPWR VPWR registers\[25\]\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_240_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21703_ _08369_ _08372_ _08062_ _08063_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__o211a_1
X_22683_ registers\[4\]\[57\] registers\[5\]\[57\] registers\[6\]\[57\] registers\[7\]\[57\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__mux4_1
X_25471_ _11015_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34669_ clknet_leaf_403_CLK _02783_ VGND VGND VPWR VPWR registers\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27210_ _11782_ registers\[37\]\[25\] _11958_ VGND VGND VPWR VPWR _11964_ sky130_fd_sc_hd__mux2_1
XFILLER_244_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24422_ net53 VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__buf_4
X_21634_ _08267_ _08304_ _08305_ _08270_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__a22o_1
X_28190_ _12480_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27141_ _11927_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__clkbuf_1
X_24353_ _10377_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
X_21565_ registers\[12\]\[25\] registers\[13\]\[25\] registers\[14\]\[25\] registers\[15\]\[25\]
+ _08173_ _08174_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__mux4_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23304_ _09708_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__buf_4
X_20516_ registers\[32\]\[62\] registers\[33\]\[62\] registers\[34\]\[62\] registers\[35\]\[62\]
+ _05108_ _05109_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__mux4_1
XFILLER_193_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24284_ registers\[57\]\[12\] _10330_ _10326_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__mux2_1
X_27072_ _11891_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21496_ _07924_ _08170_ _08171_ _07927_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__a22o_1
XFILLER_10_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26023_ _10743_ registers\[45\]\[6\] _11301_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__mux2_1
XFILLER_109_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23235_ registers\[9\]\[29\] _09751_ _09735_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__mux2_1
X_20447_ registers\[16\]\[59\] registers\[17\]\[59\] registers\[18\]\[59\] registers\[19\]\[59\]
+ _05151_ _05153_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__mux4_1
XFILLER_140_1292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_951 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23166_ _09712_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20378_ _07080_ _07083_ _06855_ _06856_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__o211a_1
XFILLER_134_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22117_ _08775_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_1208 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23097_ registers\[39\]\[3\] _09664_ _09658_ VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__mux2_1
X_27974_ _11734_ registers\[31\]\[2\] _12364_ VGND VGND VPWR VPWR _12367_ sky130_fd_sc_hd__mux2_1
XANTENNA_1219 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29713_ _13312_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__clkbuf_1
XTAP_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26925_ net27 VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__clkbuf_4
X_22048_ _08469_ _08706_ _08707_ _08472_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__a22o_1
XTAP_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29644_ registers\[20\]\[59\] _13058_ _13266_ VGND VGND VPWR VPWR _13276_ sky130_fd_sc_hd__mux2_1
XTAP_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26856_ _11752_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__clkbuf_1
XTAP_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25807_ _11194_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_235_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29575_ registers\[20\]\[26\] _12989_ _13233_ VGND VGND VPWR VPWR _13240_ sky130_fd_sc_hd__mux2_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26787_ _11710_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23999_ _10174_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_217_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28526_ _11746_ registers\[27\]\[8\] _12648_ VGND VGND VPWR VPWR _12657_ sky130_fd_sc_hd__mux2_1
X_16540_ _15037_ _15040_ _14934_ _14935_ VGND VGND VPWR VPWR _15041_ sky130_fd_sc_hd__o211a_2
X_25738_ _11156_ VGND VGND VPWR VPWR _11157_ sky130_fd_sc_hd__buf_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_216_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_243_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16471_ _14863_ _14972_ _14973_ _14867_ VGND VGND VPWR VPWR _14974_ sky130_fd_sc_hd__a22o_1
X_28457_ _12620_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25669_ registers\[48\]\[31\] _10370_ _11119_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__mux2_1
XFILLER_71_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18210_ registers\[20\]\[61\] registers\[21\]\[61\] registers\[22\]\[61\] registers\[23\]\[61\]
+ _14593_ _14595_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__mux4_1
XFILLER_223_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27408_ registers\[36\]\[55\] _10420_ _12062_ VGND VGND VPWR VPWR _12068_ sky130_fd_sc_hd__mux2_1
X_19190_ registers\[60\]\[23\] registers\[61\]\[23\] registers\[62\]\[23\] registers\[63\]\[23\]
+ _05619_ _05756_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__mux4_1
XFILLER_227_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28388_ _12584_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18141_ _14491_ _04907_ _04908_ _14501_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a22o_1
XFILLER_223_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27339_ registers\[36\]\[22\] _10351_ _12029_ VGND VGND VPWR VPWR _12032_ sky130_fd_sc_hd__mux2_1
XFILLER_12_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18072_ registers\[56\]\[57\] registers\[57\]\[57\] registers\[58\]\[57\] registers\[59\]\[57\]
+ _04751_ _04541_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__mux4_1
X_30350_ _09676_ registers\[14\]\[9\] _13638_ VGND VGND VPWR VPWR _13648_ sky130_fd_sc_hd__mux2_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29009_ registers\[24\]\[45\] _10399_ _12905_ VGND VGND VPWR VPWR _12911_ sky130_fd_sc_hd__mux2_1
X_17023_ _15341_ _15506_ _15509_ _15344_ VGND VGND VPWR VPWR _15510_ sky130_fd_sc_hd__a22o_1
XFILLER_109_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30281_ _13611_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32020_ clknet_leaf_64_CLK _00198_ VGND VGND VPWR VPWR registers\[62\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _05404_ _05718_ _05719_ _05410_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a22o_1
XANTENNA_1720 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1731 _00178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1742 _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17925_ registers\[4\]\[52\] registers\[5\]\[52\] registers\[6\]\[52\] registers\[7\]\[52\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__mux4_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33971_ clknet_leaf_349_CLK _02085_ VGND VGND VPWR VPWR registers\[37\]\[37\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1753 _07281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1764 _07843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_294_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_294_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_1775 _11753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35710_ clknet_leaf_295_CLK _03824_ VGND VGND VPWR VPWR registers\[10\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_17856_ registers\[24\]\[50\] registers\[25\]\[50\] registers\[26\]\[50\] registers\[27\]\[50\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__mux4_1
XANTENNA_1786 _14555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32922_ clknet_leaf_66_CLK _01036_ VGND VGND VPWR VPWR registers\[53\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16807_ _15295_ _15296_ _15299_ _15300_ VGND VGND VPWR VPWR _15301_ sky130_fd_sc_hd__a22o_1
XFILLER_130_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35641_ clknet_leaf_302_CLK _03755_ VGND VGND VPWR VPWR registers\[11\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_17787_ _04289_ _04564_ _04565_ _04292_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__a22o_1
X_32853_ clknet_leaf_63_CLK _00967_ VGND VGND VPWR VPWR registers\[54\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_235_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31804_ _14412_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__clkbuf_1
X_16738_ registers\[32\]\[19\] registers\[33\]\[19\] registers\[34\]\[19\] registers\[35\]\[19\]
+ _15231_ _15232_ VGND VGND VPWR VPWR _15233_ sky130_fd_sc_hd__mux4_1
X_19526_ _05127_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__buf_4
X_32784_ clknet_leaf_175_CLK _00898_ VGND VGND VPWR VPWR registers\[55\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_35572_ clknet_leaf_415_CLK _03686_ VGND VGND VPWR VPWR registers\[12\]\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34523_ clknet_leaf_1_CLK _02637_ VGND VGND VPWR VPWR registers\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_19457_ _05156_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__buf_4
X_31735_ _14376_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16669_ registers\[36\]\[17\] registers\[37\]\[17\] registers\[38\]\[17\] registers\[39\]\[17\]
+ _15164_ _15165_ VGND VGND VPWR VPWR _15166_ sky130_fd_sc_hd__mux4_1
XFILLER_223_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18408_ _05120_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31666_ registers\[63\]\[57\] net53 _14332_ VGND VGND VPWR VPWR _14340_ sky130_fd_sc_hd__mux2_1
X_34454_ clknet_leaf_87_CLK _02568_ VGND VGND VPWR VPWR registers\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_19388_ registers\[40\]\[29\] registers\[41\]\[29\] registers\[42\]\[29\] registers\[43\]\[29\]
+ _05884_ _05885_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__mux4_1
XFILLER_194_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18339_ net81 VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__buf_12
X_30617_ _13788_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__clkbuf_1
X_33405_ clknet_leaf_274_CLK _01519_ VGND VGND VPWR VPWR registers\[46\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34385_ clknet_leaf_100_CLK _02499_ VGND VGND VPWR VPWR registers\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_31597_ registers\[63\]\[24\] net17 _14299_ VGND VGND VPWR VPWR _14304_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33336_ clknet_leaf_339_CLK _01450_ VGND VGND VPWR VPWR registers\[47\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_36124_ clknet_leaf_51_CLK _04238_ VGND VGND VPWR VPWR registers\[49\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_21350_ _08026_ _08029_ _07719_ _07720_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__o211a_1
XFILLER_124_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30548_ _09773_ registers\[13\]\[39\] _13742_ VGND VGND VPWR VPWR _13752_ sky130_fd_sc_hd__mux2_1
XFILLER_129_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20301_ _06873_ _07008_ _07009_ _06878_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__a22o_1
XFILLER_162_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36055_ clknet_leaf_65_CLK _04169_ VGND VGND VPWR VPWR registers\[59\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_21281_ _07924_ _07961_ _07962_ _07927_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__a22o_1
X_33267_ clknet_leaf_364_CLK _01381_ VGND VGND VPWR VPWR registers\[48\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_30479_ _09670_ registers\[13\]\[6\] _13709_ VGND VGND VPWR VPWR _13716_ sky130_fd_sc_hd__mux2_1
XFILLER_162_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23020_ _09609_ registers\[62\]\[45\] _09599_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__mux2_1
XFILLER_239_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20232_ _05127_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__buf_4
X_32218_ clknet_leaf_292_CLK _00332_ VGND VGND VPWR VPWR registers\[9\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_35006_ clknet_leaf_188_CLK _03120_ VGND VGND VPWR VPWR registers\[21\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33198_ clknet_leaf_376_CLK _01312_ VGND VGND VPWR VPWR registers\[4\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_995 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_226_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32149_ clknet_leaf_117_CLK _00263_ VGND VGND VPWR VPWR registers\[39\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_20163_ _05093_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__buf_4
XFILLER_143_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20094_ registers\[40\]\[49\] registers\[41\]\[49\] registers\[42\]\[49\] registers\[43\]\[49\]
+ _06570_ _06571_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__mux4_1
X_24971_ _09630_ registers\[53\]\[55\] _10713_ VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__mux2_1
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_285_CLK clknet_6_56__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_285_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_26710_ _11670_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_245_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35908_ clknet_leaf_236_CLK _04022_ VGND VGND VPWR VPWR registers\[7\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_23922_ _10088_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__buf_4
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27690_ registers\[34\]\[60\] _10430_ _12150_ VGND VGND VPWR VPWR _12217_ sky130_fd_sc_hd__mux2_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26641_ _11633_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__clkbuf_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35839_ clknet_leaf_292_CLK _03953_ VGND VGND VPWR VPWR registers\[8\]\[49\] sky130_fd_sc_hd__dfxtp_1
X_23853_ _09529_ registers\[60\]\[7\] _10089_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__mux2_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_606 _05102_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _07296_ _09440_ _09441_ _07302_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__a22o_1
X_29360_ _09802_ registers\[22\]\[52\] _13124_ VGND VGND VPWR VPWR _13127_ sky130_fd_sc_hd__mux2_1
XANTENNA_617 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_246_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_232_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_628 _05122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26572_ _11585_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__clkbuf_8
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _07648_ _07684_ _07685_ _07652_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__a22o_1
X_23784_ _09596_ registers\[29\]\[39\] _10050_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__mux2_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_639 _05152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28311_ registers\[2\]\[34\] _10376_ _12539_ VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__mux2_1
X_25523_ _11042_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_241_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22735_ registers\[60\]\[59\] registers\[61\]\[59\] registers\[62\]\[59\] registers\[63\]\[59\]
+ _09227_ _07379_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__mux4_1
XFILLER_129_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29291_ _13090_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_198_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28242_ registers\[2\]\[1\] _10307_ _12506_ VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25454_ _10858_ registers\[50\]\[61\] _10936_ VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__mux2_1
X_22666_ registers\[32\]\[57\] registers\[33\]\[57\] registers\[34\]\[57\] registers\[35\]\[57\]
+ _09045_ _09046_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__mux4_1
XFILLER_197_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24405_ registers\[57\]\[51\] _10412_ _10410_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__mux2_1
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28173_ _12471_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__clkbuf_1
X_21617_ registers\[32\]\[27\] registers\[33\]\[27\] registers\[34\]\[27\] registers\[35\]\[27\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__mux4_1
X_25385_ _10789_ registers\[50\]\[28\] _10959_ VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__mux2_1
X_22597_ registers\[16\]\[54\] registers\[17\]\[54\] registers\[18\]\[54\] registers\[19\]\[54\]
+ _08965_ _08966_ VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__mux4_1
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27124_ _11918_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24336_ registers\[57\]\[29\] _10365_ _10347_ VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__mux2_1
X_21548_ _08119_ _08220_ _08221_ _08124_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__a22o_1
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27055_ _11882_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__clkbuf_1
X_24267_ net62 VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__buf_4
X_21479_ _08155_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26006_ _11298_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23218_ registers\[9\]\[24\] _09740_ _09735_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__mux2_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24198_ _10279_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23149_ _09657_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__buf_4
XANTENNA_1005 _11843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1016 _12221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1027 _12718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1038 _13139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27957_ _12357_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__clkbuf_1
XTAP_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1049 _13352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_276_CLK clknet_6_58__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_276_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17710_ _04485_ _04490_ _15974_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__o21ba_1
XFILLER_76_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26908_ _11787_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_1
X_18690_ _05440_ _05443_ _05074_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__o21ba_2
XFILLER_212_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27888_ _12321_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__clkbuf_1
XTAP_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _14562_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__buf_6
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29627_ _13267_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__clkbuf_1
X_26839_ _11740_ registers\[3\]\[5\] _11730_ VGND VGND VPWR VPWR _11741_ sky130_fd_sc_hd__mux2_1
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17572_ registers\[4\]\[42\] registers\[5\]\[42\] registers\[6\]\[42\] registers\[7\]\[42\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__mux4_1
X_29558_ registers\[20\]\[18\] _12972_ _13222_ VGND VGND VPWR VPWR _13231_ sky130_fd_sc_hd__mux2_1
XFILLER_223_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19311_ registers\[20\]\[26\] registers\[21\]\[26\] registers\[22\]\[26\] registers\[23\]\[26\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__mux4_1
X_28509_ _12647_ VGND VGND VPWR VPWR _12648_ sky130_fd_sc_hd__buf_4
XFILLER_204_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16523_ _14952_ _15023_ _15024_ _14957_ VGND VGND VPWR VPWR _15025_ sky130_fd_sc_hd__a22o_1
XFILLER_189_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_232_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29489_ _13194_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31520_ _14263_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19242_ _05844_ _05979_ _05980_ _05849_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__a22o_1
XFILLER_220_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16454_ _14952_ _14953_ _14956_ _14957_ VGND VGND VPWR VPWR _14958_ sky130_fd_sc_hd__a22o_1
XFILLER_91_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31451_ _09697_ registers\[6\]\[19\] _14217_ VGND VGND VPWR VPWR _14227_ sky130_fd_sc_hd__mux2_1
X_19173_ _05152_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__clkbuf_4
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16385_ registers\[32\]\[9\] registers\[33\]\[9\] registers\[34\]\[9\] registers\[35\]\[9\]
+ _14888_ _14889_ VGND VGND VPWR VPWR _14890_ sky130_fd_sc_hd__mux4_1
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_200_CLK clknet_6_51__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_200_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18124_ _04892_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_2
X_30402_ _13675_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__clkbuf_1
X_34170_ clknet_leaf_281_CLK _02284_ VGND VGND VPWR VPWR registers\[34\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_31382_ registers\[7\]\[50\] net46 _14190_ VGND VGND VPWR VPWR _14191_ sky130_fd_sc_hd__mux2_1
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33121_ clknet_leaf_42_CLK _01235_ VGND VGND VPWR VPWR registers\[50\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_18055_ _04822_ _04825_ _04630_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__o21ba_1
X_30333_ _13639_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ _14592_ VGND VGND VPWR VPWR _15494_ sky130_fd_sc_hd__buf_4
X_33052_ clknet_leaf_51_CLK _01166_ VGND VGND VPWR VPWR registers\[51\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_30264_ _13602_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32003_ clknet_leaf_28_CLK _00176_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30195_ _13565_ VGND VGND VPWR VPWR _13566_ sky130_fd_sc_hd__buf_4
XFILLER_99_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18957_ registers\[28\]\[16\] registers\[29\]\[16\] registers\[30\]\[16\] registers\[31\]\[16\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__mux4_1
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_230_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_267_CLK clknet_6_57__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_267_CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_1550 _11300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1561 _11585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ _14539_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__buf_4
XANTENNA_1572 _12972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1583 _14276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33954_ clknet_leaf_47_CLK _02068_ VGND VGND VPWR VPWR registers\[37\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_18888_ registers\[20\]\[14\] registers\[21\]\[14\] registers\[22\]\[14\] registers\[23\]\[14\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__mux4_1
XFILLER_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1594 _14539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32905_ clknet_leaf_177_CLK _01019_ VGND VGND VPWR VPWR registers\[54\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_17839_ registers\[60\]\[50\] registers\[61\]\[50\] registers\[62\]\[50\] registers\[63\]\[50\]
+ _04412_ _04549_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__mux4_1
X_33885_ clknet_leaf_22_CLK _01999_ VGND VGND VPWR VPWR registers\[38\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_20850_ registers\[60\]\[5\] registers\[61\]\[5\] registers\[62\]\[5\] registers\[63\]\[5\]
+ _07512_ _07329_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__mux4_1
X_35624_ clknet_leaf_460_CLK _03738_ VGND VGND VPWR VPWR registers\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_32836_ clknet_leaf_200_CLK _00950_ VGND VGND VPWR VPWR registers\[55\]\[54\] sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19509_ registers\[48\]\[32\] registers\[49\]\[32\] registers\[50\]\[32\] registers\[51\]\[32\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux4_1
X_20781_ registers\[56\]\[3\] registers\[57\]\[3\] registers\[58\]\[3\] registers\[59\]\[3\]
+ _07315_ _07317_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__mux4_1
X_35555_ clknet_leaf_469_CLK _03669_ VGND VGND VPWR VPWR registers\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32767_ clknet_leaf_268_CLK _00881_ VGND VGND VPWR VPWR registers\[56\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34506_ clknet_leaf_153_CLK _02620_ VGND VGND VPWR VPWR registers\[2\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_223_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22520_ _09163_ _09166_ _09091_ _09092_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__o211a_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31718_ _14367_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32698_ clknet_leaf_285_CLK _00812_ VGND VGND VPWR VPWR registers\[57\]\[44\] sky130_fd_sc_hd__dfxtp_1
X_35486_ clknet_leaf_483_CLK _03600_ VGND VGND VPWR VPWR registers\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34437_ clknet_leaf_213_CLK _02551_ VGND VGND VPWR VPWR registers\[30\]\[55\] sky130_fd_sc_hd__dfxtp_1
X_22451_ registers\[4\]\[50\] registers\[5\]\[50\] registers\[6\]\[50\] registers\[7\]\[50\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__mux4_1
X_31649_ registers\[63\]\[49\] net44 _14321_ VGND VGND VPWR VPWR _14331_ sky130_fd_sc_hd__mux2_1
XFILLER_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21402_ registers\[28\]\[20\] registers\[29\]\[20\] registers\[30\]\[20\] registers\[31\]\[20\]
+ _07806_ _07807_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__mux4_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25170_ _10851_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__clkbuf_1
X_22382_ registers\[4\]\[48\] registers\[5\]\[48\] registers\[6\]\[48\] registers\[7\]\[48\]
+ _09031_ _09032_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__mux4_1
X_34368_ clknet_leaf_199_CLK _02482_ VGND VGND VPWR VPWR registers\[31\]\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36107_ clknet_leaf_164_CLK _04221_ VGND VGND VPWR VPWR registers\[59\]\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24121_ _09525_ registers\[58\]\[5\] _10233_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__mux2_1
X_21333_ _07982_ _07997_ _08006_ _08013_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__or4_2
X_33319_ clknet_leaf_60_CLK _01433_ VGND VGND VPWR VPWR registers\[47\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_34299_ clknet_leaf_279_CLK _02413_ VGND VGND VPWR VPWR registers\[32\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36038_ clknet_leaf_194_CLK _04152_ VGND VGND VPWR VPWR registers\[63\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_24052_ _09592_ registers\[5\]\[37\] _10194_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__mux2_1
X_21264_ registers\[32\]\[17\] registers\[33\]\[17\] registers\[34\]\[17\] registers\[35\]\[17\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__mux4_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20215_ registers\[48\]\[52\] registers\[49\]\[52\] registers\[50\]\[52\] registers\[51\]\[52\]
+ _06779_ _06780_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__mux4_1
X_23003_ net35 VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__clkbuf_4
Xmax_cap282 _12860_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_12
XFILLER_176_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28860_ _12832_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__clkbuf_1
X_21195_ _07776_ _07877_ _07878_ _07781_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__a22o_1
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_235_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27811_ registers\[33\]\[53\] _10416_ _12277_ VGND VGND VPWR VPWR _12281_ sky130_fd_sc_hd__mux2_1
X_20146_ _05120_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__buf_6
X_28791_ _12796_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_258_CLK clknet_6_62__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_258_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ registers\[33\]\[20\] _10346_ _12244_ VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__mux2_1
X_20077_ registers\[0\]\[48\] registers\[1\]\[48\] registers\[2\]\[48\] registers\[3\]\[48\]
+ _06516_ _06517_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__mux4_1
X_24954_ _09613_ registers\[53\]\[47\] _10702_ VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__mux2_1
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_840 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_6_27__f_CLK clknet_5_13_0_CLK VGND VGND VPWR VPWR clknet_6_27__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _10124_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27673_ _12208_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__clkbuf_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24885_ _09544_ registers\[53\]\[14\] _10669_ VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__mux2_1
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_248_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_233_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29412_ _13154_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__clkbuf_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26624_ _11624_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__clkbuf_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _09941_ net83 _09512_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__or3b_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_908 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_436 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29343_ _09784_ registers\[22\]\[44\] _13113_ VGND VGND VPWR VPWR _13118_ sky130_fd_sc_hd__mux2_1
XANTENNA_447 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26555_ _11588_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_458 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23767_ _10051_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20979_ _07666_ _07669_ _07399_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__o21ba_1
XANTENNA_469 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_430_CLK clknet_6_15__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_430_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25506_ _11033_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__clkbuf_1
X_22718_ _09104_ _09357_ _09358_ _09107_ VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__a22o_1
XFILLER_213_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29274_ _09681_ registers\[22\]\[11\] _13080_ VGND VGND VPWR VPWR _13082_ sky130_fd_sc_hd__mux2_1
XFILLER_201_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26486_ _11551_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__clkbuf_1
X_23698_ _09649_ _09650_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__nand2_2
XFILLER_158_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28225_ _12498_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__clkbuf_1
X_25437_ _10995_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22649_ registers\[8\]\[56\] registers\[9\]\[56\] registers\[10\]\[56\] registers\[11\]\[56\]
+ _07288_ _07290_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__mux4_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16170_ _14601_ _14680_ _14681_ _14611_ VGND VGND VPWR VPWR _14682_ sky130_fd_sc_hd__a22o_1
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28156_ _12462_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25368_ _10936_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__buf_4
XFILLER_220_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27107_ _11813_ registers\[38\]\[40\] _11909_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__mux2_1
X_24319_ _10354_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
X_28087_ _11847_ registers\[31\]\[56\] _12419_ VGND VGND VPWR VPWR _12426_ sky130_fd_sc_hd__mux2_1
X_25299_ _10922_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__clkbuf_1
X_27038_ _11873_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19860_ _06575_ _06580_ _06504_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__o21ba_1
X_18811_ _05345_ _05560_ _05561_ _05348_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__a22o_1
XTAP_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput94 net94 VGND VGND VPWR VPWR D1[13] sky130_fd_sc_hd__buf_2
X_19791_ _06508_ _06511_ _06512_ _06513_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__o211a_1
XTAP_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28989_ _12900_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_249_CLK clknet_6_63__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_249_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18742_ _05490_ _05493_ _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__o21ba_1
XFILLER_231_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18673_ registers\[24\]\[8\] registers\[25\]\[8\] registers\[26\]\[8\] registers\[27\]\[8\]
+ _05288_ _05289_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__mux4_1
X_30951_ registers\[10\]\[38\] _13014_ _13955_ VGND VGND VPWR VPWR _13964_ sky130_fd_sc_hd__mux2_1
XFILLER_97_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _04403_ _04406_ _15955_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__o21ba_1
X_33670_ clknet_leaf_248_CLK _01784_ VGND VGND VPWR VPWR registers\[42\]\[56\] sky130_fd_sc_hd__dfxtp_1
X_30882_ registers\[10\]\[5\] _12945_ _13922_ VGND VGND VPWR VPWR _13928_ sky130_fd_sc_hd__mux2_1
XFILLER_40_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _14539_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__clkbuf_4
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32621_ clknet_leaf_372_CLK _00735_ VGND VGND VPWR VPWR registers\[58\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16506_ registers\[52\]\[12\] registers\[53\]\[12\] registers\[54\]\[12\] registers\[55\]\[12\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _15008_ sky130_fd_sc_hd__mux4_1
XANTENNA_970 _11011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_421_CLK clknet_6_36__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_421_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_35340_ clknet_leaf_148_CLK _03454_ VGND VGND VPWR VPWR registers\[16\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_981 _11300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_32552_ clknet_leaf_401_CLK _00666_ VGND VGND VPWR VPWR registers\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_992 _11738_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17486_ registers\[60\]\[40\] registers\[61\]\[40\] registers\[62\]\[40\] registers\[63\]\[40\]
+ _15756_ _15893_ VGND VGND VPWR VPWR _15960_ sky130_fd_sc_hd__mux4_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31503_ _14254_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_220_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16437_ _14796_ _14937_ _14940_ _14799_ VGND VGND VPWR VPWR _14941_ sky130_fd_sc_hd__a22o_1
X_19225_ registers\[52\]\[24\] registers\[53\]\[24\] registers\[54\]\[24\] registers\[55\]\[24\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__mux4_1
X_35271_ clknet_leaf_153_CLK _03385_ VGND VGND VPWR VPWR registers\[17\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32483_ clknet_leaf_445_CLK _00597_ VGND VGND VPWR VPWR registers\[60\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31434_ _14218_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__clkbuf_1
X_34222_ clknet_leaf_352_CLK _02336_ VGND VGND VPWR VPWR registers\[33\]\[32\] sky130_fd_sc_hd__dfxtp_1
X_19156_ registers\[48\]\[22\] registers\[49\]\[22\] registers\[50\]\[22\] registers\[51\]\[22\]
+ _05750_ _05751_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__mux4_1
X_16368_ _14576_ VGND VGND VPWR VPWR _14874_ sky130_fd_sc_hd__buf_6
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18107_ _14600_ _04874_ _04875_ _14610_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__a22o_1
XFILLER_30_1129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34153_ clknet_leaf_431_CLK _02267_ VGND VGND VPWR VPWR registers\[34\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31365_ registers\[7\]\[42\] net37 _14179_ VGND VGND VPWR VPWR _14182_ sky130_fd_sc_hd__mux2_1
X_19087_ _05111_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__buf_6
X_16299_ registers\[24\]\[6\] registers\[25\]\[6\] registers\[26\]\[6\] registers\[27\]\[6\]
+ _14739_ _14740_ VGND VGND VPWR VPWR _14807_ sky130_fd_sc_hd__mux4_1
XFILLER_69_1328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30316_ _13629_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__clkbuf_1
X_18038_ registers\[44\]\[56\] registers\[45\]\[56\] registers\[46\]\[56\] registers\[47\]\[56\]
+ _04606_ _04607_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__mux4_1
X_33104_ clknet_leaf_75_CLK _01218_ VGND VGND VPWR VPWR registers\[50\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_34084_ clknet_leaf_56_CLK _02198_ VGND VGND VPWR VPWR registers\[35\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_31296_ _14145_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_488_CLK clknet_6_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_488_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_33035_ clknet_leaf_165_CLK _01149_ VGND VGND VPWR VPWR registers\[52\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_30247_ _13593_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_236_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20000_ _05039_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__buf_4
X_30178_ registers\[16\]\[56\] _13052_ _13550_ VGND VGND VPWR VPWR _13557_ sky130_fd_sc_hd__mux2_1
X_19989_ _06576_ _06704_ _06705_ _06579_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__a22o_1
XFILLER_143_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34986_ clknet_leaf_453_CLK _03100_ VGND VGND VPWR VPWR registers\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1380 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_239_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1391 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33937_ clknet_leaf_134_CLK _02051_ VGND VGND VPWR VPWR registers\[37\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21951_ _08610_ _08611_ _08612_ _08613_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__a22o_1
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ registers\[16\]\[6\] registers\[17\]\[6\] registers\[18\]\[6\] registers\[19\]\[6\]
+ _07593_ _07594_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__mux4_1
X_24670_ _09601_ registers\[55\]\[41\] _10558_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__mux2_1
X_33868_ clknet_leaf_148_CLK _01982_ VGND VGND VPWR VPWR registers\[3\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_21882_ registers\[0\]\[34\] registers\[1\]\[34\] registers\[2\]\[34\] registers\[3\]\[34\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__mux4_1
XFILLER_55_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35607_ clknet_leaf_87_CLK _03721_ VGND VGND VPWR VPWR registers\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ registers\[61\]\[27\] _09747_ _09965_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__mux2_1
X_20833_ _07373_ _07526_ _07527_ _07383_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__a22o_1
X_32819_ clknet_leaf_355_CLK _00933_ VGND VGND VPWR VPWR registers\[55\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_208_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33799_ clknet_leaf_243_CLK _01913_ VGND VGND VPWR VPWR registers\[40\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_230_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_412_CLK clknet_6_35__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_412_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26340_ _11474_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__clkbuf_1
X_23552_ _09935_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35538_ clknet_leaf_107_CLK _03652_ VGND VGND VPWR VPWR registers\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20764_ registers\[16\]\[2\] registers\[17\]\[2\] registers\[18\]\[2\] registers\[19\]\[2\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__mux4_1
XFILLER_11_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22503_ _07281_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__buf_6
XFILLER_195_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26271_ _10856_ registers\[44\]\[60\] _11371_ VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__mux2_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35469_ clknet_leaf_133_CLK _03583_ VGND VGND VPWR VPWR registers\[14\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_20695_ registers\[20\]\[0\] registers\[21\]\[0\] registers\[22\]\[0\] registers\[23\]\[0\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__mux4_1
X_23483_ _09899_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28010_ _12385_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25222_ _10762_ registers\[51\]\[15\] _10876_ VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__mux2_1
X_22434_ _07309_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__buf_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_195_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_17_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_17_0_CLK sky130_fd_sc_hd__clkbuf_8
X_25153_ net48 VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_104_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22365_ _07328_ VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_191_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24104_ _09644_ registers\[5\]\[62\] _10160_ VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__mux2_1
XFILLER_124_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21316_ _07990_ _07996_ _07719_ _07720_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__o211a_1
X_22296_ _07333_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__clkbuf_4
XFILLER_164_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25084_ net24 VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__buf_4
X_29961_ registers\[17\]\[17\] _12970_ _13435_ VGND VGND VPWR VPWR _13443_ sky130_fd_sc_hd__mux2_1
XFILLER_190_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_479_CLK clknet_6_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_479_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28912_ _12859_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__clkbuf_1
X_21247_ registers\[12\]\[16\] registers\[13\]\[16\] registers\[14\]\[16\] registers\[15\]\[16\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__mux4_1
X_24035_ _09575_ registers\[5\]\[29\] _10183_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__mux2_1
XFILLER_85_1152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29892_ _13406_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21178_ registers\[12\]\[14\] registers\[13\]\[14\] registers\[14\]\[14\] registers\[15\]\[14\]
+ _07830_ _07831_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__mux4_1
X_28843_ _11792_ registers\[25\]\[30\] _12823_ VGND VGND VPWR VPWR _12824_ sky130_fd_sc_hd__mux2_1
XFILLER_137_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20129_ _05095_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__buf_4
XFILLER_77_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28774_ _11859_ registers\[26\]\[62\] _12718_ VGND VGND VPWR VPWR _12787_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25986_ _11288_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27725_ registers\[33\]\[12\] _10330_ _12233_ VGND VGND VPWR VPWR _12236_ sky130_fd_sc_hd__mux2_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24937_ _09596_ registers\[53\]\[39\] _10691_ VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__mux2_1
XFILLER_213_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27656_ _12199_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24868_ _09527_ registers\[53\]\[6\] _10658_ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__mux2_1
XANTENNA_200 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26607_ _11615_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__clkbuf_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23819_ _10078_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_233 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27587_ _12163_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__clkbuf_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_255 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24799_ _10628_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_266 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_403_CLK clknet_6_33__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_403_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_277 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17340_ _15541_ _15816_ _15817_ _15547_ VGND VGND VPWR VPWR _15818_ sky130_fd_sc_hd__a22o_1
X_29326_ _09766_ registers\[22\]\[36\] _13102_ VGND VGND VPWR VPWR _13109_ sky130_fd_sc_hd__mux2_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26538_ _11578_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_288 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_299 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29257_ _09664_ registers\[22\]\[3\] _13069_ VGND VGND VPWR VPWR _13073_ sky130_fd_sc_hd__mux2_1
X_17271_ _15747_ _15750_ _15612_ VGND VGND VPWR VPWR _15751_ sky130_fd_sc_hd__o21ba_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26469_ _11542_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19010_ _05088_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__clkbuf_4
X_16222_ registers\[8\]\[4\] registers\[9\]\[4\] registers\[10\]\[4\] registers\[11\]\[4\]
+ _14559_ _14560_ VGND VGND VPWR VPWR _14732_ sky130_fd_sc_hd__mux4_1
X_28208_ _12489_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29188_ net39 VGND VGND VPWR VPWR _13027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16153_ registers\[52\]\[2\] registers\[53\]\[2\] registers\[54\]\[2\] registers\[55\]\[2\]
+ _14547_ _14549_ VGND VGND VPWR VPWR _14665_ sky130_fd_sc_hd__mux4_1
X_28139_ _12453_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31150_ registers\[8\]\[4\] net45 _14064_ VGND VGND VPWR VPWR _14069_ sky130_fd_sc_hd__mux2_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16084_ _14597_ VGND VGND VPWR VPWR _14598_ sky130_fd_sc_hd__buf_4
XFILLER_6_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1077 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30101_ _13516_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__clkbuf_1
X_19912_ registers\[28\]\[43\] registers\[29\]\[43\] registers\[30\]\[43\] registers\[31\]\[43\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__mux4_1
XFILLER_218_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_31081_ _14032_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1052 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30032_ _13480_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__clkbuf_1
X_19843_ registers\[20\]\[41\] registers\[21\]\[41\] registers\[22\]\[41\] registers\[23\]\[41\]
+ _06532_ _06533_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__mux4_1
XFILLER_64_1247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34840_ clknet_leaf_2_CLK _02954_ VGND VGND VPWR VPWR registers\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19774_ registers\[32\]\[40\] registers\[33\]\[40\] registers\[34\]\[40\] registers\[35\]\[40\]
+ _06466_ _06467_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__mux4_1
X_16986_ registers\[48\]\[26\] registers\[49\]\[26\] registers\[50\]\[26\] registers\[51\]\[26\]
+ _15201_ _15202_ VGND VGND VPWR VPWR _15474_ sky130_fd_sc_hd__mux4_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_231_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18725_ registers\[48\]\[10\] registers\[49\]\[10\] registers\[50\]\[10\] registers\[51\]\[10\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__mux4_1
XFILLER_231_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34771_ clknet_leaf_80_CLK _02885_ VGND VGND VPWR VPWR registers\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31983_ clknet_leaf_21_CLK _00154_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_237_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33722_ clknet_leaf_279_CLK _01836_ VGND VGND VPWR VPWR registers\[41\]\[44\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_6_10__f_CLK clknet_5_5_0_CLK VGND VGND VPWR VPWR clknet_6_10__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_18656_ _05404_ _05406_ _05409_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a22o_1
X_30934_ _13921_ VGND VGND VPWR VPWR _13955_ sky130_fd_sc_hd__buf_4
XFILLER_188_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17607_ _15830_ _04389_ _04390_ _15833_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__a22o_1
X_30865_ _13918_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_33653_ clknet_leaf_343_CLK _01767_ VGND VGND VPWR VPWR registers\[42\]\[39\] sky130_fd_sc_hd__dfxtp_1
X_18587_ _05338_ _05343_ _05103_ _05105_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__o211a_1
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_233_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_32604_ clknet_leaf_37_CLK _00718_ VGND VGND VPWR VPWR registers\[58\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_17538_ _04320_ _04323_ _15974_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__o21ba_1
X_30796_ _13882_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__clkbuf_1
X_33584_ clknet_leaf_347_CLK _01698_ VGND VGND VPWR VPWR registers\[43\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35323_ clknet_leaf_186_CLK _03437_ VGND VGND VPWR VPWR registers\[16\]\[45\] sky130_fd_sc_hd__dfxtp_1
X_32535_ clknet_leaf_83_CLK _00649_ VGND VGND VPWR VPWR registers\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_17469_ _15638_ _15942_ _15943_ _15643_ VGND VGND VPWR VPWR _15944_ sky130_fd_sc_hd__a22o_1
XFILLER_203_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19208_ _05844_ _05946_ _05947_ _05849_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a22o_1
X_20480_ registers\[20\]\[60\] registers\[21\]\[60\] registers\[22\]\[60\] registers\[23\]\[60\]
+ _05142_ _05144_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__mux4_1
XFILLER_165_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35254_ clknet_leaf_310_CLK _03368_ VGND VGND VPWR VPWR registers\[17\]\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32466_ clknet_leaf_181_CLK _00580_ VGND VGND VPWR VPWR registers\[60\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34205_ clknet_leaf_22_CLK _02319_ VGND VGND VPWR VPWR registers\[33\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_31417_ _14209_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__clkbuf_1
X_19139_ _05877_ _05880_ _05851_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__o21ba_1
X_32397_ clknet_leaf_167_CLK _00511_ VGND VGND VPWR VPWR registers\[61\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_35185_ clknet_leaf_395_CLK _03299_ VGND VGND VPWR VPWR registers\[18\]\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22150_ _07281_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__clkbuf_4
X_34136_ clknet_leaf_86_CLK _02250_ VGND VGND VPWR VPWR registers\[34\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_31348_ registers\[7\]\[34\] net28 _14168_ VGND VGND VPWR VPWR _14173_ sky130_fd_sc_hd__mux2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21101_ _07782_ _07787_ _07711_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__o21ba_1
X_22081_ _07309_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__buf_2
XTAP_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34067_ clknet_leaf_120_CLK _02181_ VGND VGND VPWR VPWR registers\[35\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_31279_ registers\[7\]\[1\] net12 _14135_ VGND VGND VPWR VPWR _14137_ sky130_fd_sc_hd__mux2_1
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21032_ _07715_ _07718_ _07719_ _07720_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__o211a_1
X_33018_ clknet_leaf_285_CLK _01132_ VGND VGND VPWR VPWR registers\[52\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_236_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25840_ _11211_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_247_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25771_ _11175_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22983_ _09584_ registers\[62\]\[33\] _09578_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__mux2_1
X_34969_ clknet_leaf_3_CLK _03083_ VGND VGND VPWR VPWR registers\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27510_ _12121_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__clkbuf_1
X_24722_ _10588_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__clkbuf_1
X_28490_ _11845_ registers\[28\]\[55\] _12632_ VGND VGND VPWR VPWR _12638_ sky130_fd_sc_hd__mux2_1
X_21934_ registers\[44\]\[36\] registers\[45\]\[36\] registers\[46\]\[36\] registers\[47\]\[36\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__mux4_1
XFILLER_103_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_874 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27441_ _12085_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24653_ _09584_ registers\[55\]\[33\] _10547_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__mux2_1
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ registers\[40\]\[34\] registers\[41\]\[34\] registers\[42\]\[34\] registers\[43\]\[34\]
+ _08463_ _08464_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__mux4_1
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ registers\[61\]\[19\] _09697_ _09954_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__mux2_1
X_20816_ _07313_ _07509_ _07510_ _07322_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__a22o_1
X_27372_ registers\[36\]\[38\] _10384_ _12040_ VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__mux2_1
X_24584_ _09510_ registers\[55\]\[0\] _10514_ VGND VGND VPWR VPWR _10515_ sky130_fd_sc_hd__mux2_1
XFILLER_93_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21796_ _07278_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__buf_4
XFILLER_230_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29111_ registers\[23\]\[19\] _12974_ _12956_ VGND VGND VPWR VPWR _12975_ sky130_fd_sc_hd__mux2_1
XFILLER_11_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_0_0_CLK clknet_2_0_0_CLK VGND VGND VPWR VPWR clknet_5_0_0_CLK sky130_fd_sc_hd__clkbuf_8
X_26323_ _10772_ registers\[43\]\[20\] _11465_ VGND VGND VPWR VPWR _11466_ sky130_fd_sc_hd__mux2_1
X_23535_ _09622_ registers\[19\]\[51\] _09925_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__mux2_1
X_20747_ _07440_ _07441_ _07442_ _07443_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__a22o_1
X_29042_ registers\[24\]\[61\] _10432_ _12860_ VGND VGND VPWR VPWR _12928_ sky130_fd_sc_hd__mux2_1
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26254_ _11429_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23466_ _09890_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__clkbuf_1
X_20678_ _07314_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__buf_12
XFILLER_17_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25205_ _10745_ registers\[51\]\[7\] _10865_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__mux2_1
X_22417_ registers\[24\]\[49\] registers\[25\]\[49\] registers\[26\]\[49\] registers\[27\]\[49\]
+ _08896_ _08897_ VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__mux4_1
X_26185_ _10770_ registers\[44\]\[19\] _11383_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__mux2_1
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23397_ registers\[39\]\[51\] _09800_ _09851_ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__mux2_1
X_25136_ _10828_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__clkbuf_1
X_22348_ registers\[28\]\[47\] registers\[29\]\[47\] registers\[30\]\[47\] registers\[31\]\[47\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__mux4_1
XFILLER_174_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29944_ registers\[17\]\[9\] _12953_ _13424_ VGND VGND VPWR VPWR _13434_ sky130_fd_sc_hd__mux2_1
X_25067_ _10781_ registers\[52\]\[24\] _10773_ VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__mux2_1
X_22279_ registers\[20\]\[45\] registers\[21\]\[45\] registers\[22\]\[45\] registers\[23\]\[45\]
+ _08768_ _08769_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__mux4_1
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24018_ _10184_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_239_906 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29875_ registers\[18\]\[40\] _13018_ _13397_ VGND VGND VPWR VPWR _13398_ sky130_fd_sc_hd__mux2_1
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28826_ _11776_ registers\[25\]\[22\] _12812_ VGND VGND VPWR VPWR _12815_ sky130_fd_sc_hd__mux2_1
X_16840_ _15311_ _15318_ _15325_ _15332_ VGND VGND VPWR VPWR _15333_ sky130_fd_sc_hd__or4_4
XFILLER_120_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16771_ _14548_ VGND VGND VPWR VPWR _15265_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28757_ _12778_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25969_ _11279_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_219_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18510_ registers\[36\]\[4\] registers\[37\]\[4\] registers\[38\]\[4\] registers\[39\]\[4\]
+ _05170_ _05171_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__mux4_1
XFILLER_219_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27708_ registers\[33\]\[4\] _10313_ _12222_ VGND VGND VPWR VPWR _12227_ sky130_fd_sc_hd__mux2_1
XFILLER_189_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19490_ registers\[20\]\[31\] registers\[21\]\[31\] registers\[22\]\[31\] registers\[23\]\[31\]
+ _06189_ _06190_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__mux4_1
XFILLER_46_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28688_ _12742_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__clkbuf_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18441_ _05116_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__clkbuf_8
XFILLER_111_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_896 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27639_ _12190_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__clkbuf_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _05118_ _05132_ _05134_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__o21ba_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30650_ registers\[12\]\[23\] _12983_ _13802_ VGND VGND VPWR VPWR _13806_ sky130_fd_sc_hd__mux2_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ registers\[16\]\[35\] registers\[17\]\[35\] registers\[18\]\[35\] registers\[19\]\[35\]
+ _15494_ _15495_ VGND VGND VPWR VPWR _15802_ sky130_fd_sc_hd__mux4_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29309_ _09749_ registers\[22\]\[28\] _13091_ VGND VGND VPWR VPWR _13100_ sky130_fd_sc_hd__mux2_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30581_ _13769_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__clkbuf_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32320_ clknet_leaf_221_CLK _00434_ VGND VGND VPWR VPWR registers\[19\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_17254_ _15487_ _15733_ _15734_ _15490_ VGND VGND VPWR VPWR _15735_ sky130_fd_sc_hd__a22o_1
XFILLER_105_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16205_ _14715_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32251_ clknet_leaf_282_CLK _00365_ VGND VGND VPWR VPWR registers\[39\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17185_ _15664_ _15667_ _15631_ VGND VGND VPWR VPWR _15668_ sky130_fd_sc_hd__o21ba_1
X_31202_ registers\[8\]\[29\] net22 _14086_ VGND VGND VPWR VPWR _14096_ sky130_fd_sc_hd__mux2_1
X_16136_ _14490_ VGND VGND VPWR VPWR _14648_ sky130_fd_sc_hd__buf_4
X_32182_ clknet_leaf_440_CLK _00296_ VGND VGND VPWR VPWR registers\[39\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31133_ _14059_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16067_ _14515_ VGND VGND VPWR VPWR _14581_ sky130_fd_sc_hd__buf_12
XFILLER_9_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1011 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31064_ _14023_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__clkbuf_1
X_35941_ clknet_leaf_464_CLK _04055_ VGND VGND VPWR VPWR registers\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30015_ _13471_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__clkbuf_1
X_19826_ registers\[48\]\[41\] registers\[49\]\[41\] registers\[50\]\[41\] registers\[51\]\[41\]
+ _06436_ _06437_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__mux4_1
X_35872_ clknet_leaf_468_CLK _03986_ VGND VGND VPWR VPWR registers\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_229_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34823_ clknet_leaf_219_CLK _02937_ VGND VGND VPWR VPWR registers\[24\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19757_ registers\[8\]\[39\] registers\[9\]\[39\] registers\[10\]\[39\] registers\[11\]\[39\]
+ _06341_ _06342_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__mux4_1
X_16969_ registers\[24\]\[25\] registers\[25\]\[25\] registers\[26\]\[25\] registers\[27\]\[25\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15458_ sky130_fd_sc_hd__mux4_1
X_18708_ registers\[28\]\[9\] registers\[29\]\[9\] registers\[30\]\[9\] registers\[31\]\[9\]
+ _05227_ _05228_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__mux4_1
X_34754_ clknet_leaf_224_CLK _02868_ VGND VGND VPWR VPWR registers\[25\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_31966_ clknet_leaf_4_CLK _00135_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
X_19688_ registers\[12\]\[37\] registers\[13\]\[37\] registers\[14\]\[37\] registers\[15\]\[37\]
+ _06280_ _06281_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux4_1
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33705_ clknet_leaf_428_CLK _01819_ VGND VGND VPWR VPWR registers\[41\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_213_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18639_ _05391_ _05394_ _05163_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__o21ba_1
X_30917_ _13946_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34685_ clknet_leaf_183_CLK _02799_ VGND VGND VPWR VPWR registers\[26\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31897_ _14461_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_212_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21650_ _08119_ _08319_ _08320_ _08124_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__a22o_1
X_33636_ clknet_leaf_56_CLK _01750_ VGND VGND VPWR VPWR registers\[42\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_30848_ _09804_ registers\[11\]\[53\] _13906_ VGND VGND VPWR VPWR _13910_ sky130_fd_sc_hd__mux2_1
XFILLER_127_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_244_1465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_221_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20601_ net74 net73 VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__nor2b_4
X_21581_ registers\[44\]\[26\] registers\[45\]\[26\] registers\[46\]\[26\] registers\[47\]\[26\]
+ _08049_ _08050_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__mux4_1
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33567_ clknet_leaf_33_CLK _01681_ VGND VGND VPWR VPWR registers\[43\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_30779_ _09699_ registers\[11\]\[20\] _13873_ VGND VGND VPWR VPWR _13874_ sky130_fd_sc_hd__mux2_1
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23320_ registers\[9\]\[55\] _09808_ _09798_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__mux2_1
XFILLER_221_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35306_ clknet_leaf_406_CLK _03420_ VGND VGND VPWR VPWR registers\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20532_ registers\[12\]\[62\] registers\[13\]\[62\] registers\[14\]\[62\] registers\[15\]\[62\]
+ _06966_ _06967_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__mux4_1
X_32518_ clknet_leaf_195_CLK _00632_ VGND VGND VPWR VPWR registers\[60\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33498_ clknet_leaf_31_CLK _01612_ VGND VGND VPWR VPWR registers\[44\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20463_ registers\[48\]\[60\] registers\[49\]\[60\] registers\[50\]\[60\] registers\[51\]\[60\]
+ _05091_ _05156_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__mux4_1
X_23251_ registers\[9\]\[34\] _09762_ _09754_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__mux2_1
X_35237_ clknet_leaf_448_CLK _03351_ VGND VGND VPWR VPWR registers\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_32449_ clknet_leaf_199_CLK _00563_ VGND VGND VPWR VPWR registers\[29\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22202_ _08610_ _08856_ _08857_ _08613_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__a22o_1
XFILLER_134_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20394_ _07099_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__buf_4
X_23182_ registers\[9\]\[9\] _09676_ _09709_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__mux2_1
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35168_ clknet_leaf_1_CLK _03282_ VGND VGND VPWR VPWR registers\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34119_ clknet_leaf_244_CLK _02233_ VGND VGND VPWR VPWR registers\[35\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22133_ registers\[0\]\[41\] registers\[1\]\[41\] registers\[2\]\[41\] registers\[3\]\[41\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__mux4_1
X_27990_ _12363_ VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__buf_4
X_35099_ clknet_leaf_479_CLK _03213_ VGND VGND VPWR VPWR registers\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xoutput240 net240 VGND VGND VPWR VPWR D3[2] sky130_fd_sc_hd__buf_2
XTAP_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput251 net251 VGND VGND VPWR VPWR D3[3] sky130_fd_sc_hd__buf_2
XTAP_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput262 net262 VGND VGND VPWR VPWR D3[4] sky130_fd_sc_hd__buf_2
XTAP_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26941_ _11809_ registers\[3\]\[38\] _11793_ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__mux2_1
XTAP_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput273 net273 VGND VGND VPWR VPWR D3[5] sky130_fd_sc_hd__buf_2
X_22064_ registers\[24\]\[39\] registers\[25\]\[39\] registers\[26\]\[39\] registers\[27\]\[39\]
+ _08553_ _08554_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__mux4_1
XFILLER_160_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21015_ registers\[32\]\[10\] registers\[33\]\[10\] registers\[34\]\[10\] registers\[35\]\[10\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__mux4_1
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29660_ registers\[1\]\[2\] _12939_ _13282_ VGND VGND VPWR VPWR _13285_ sky130_fd_sc_hd__mux2_1
XTAP_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26872_ net8 VGND VGND VPWR VPWR _11763_ sky130_fd_sc_hd__buf_4
XTAP_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28611_ _12701_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__clkbuf_1
X_25823_ _11202_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
X_29591_ _13248_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25754_ _11166_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_228_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28542_ _12665_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__clkbuf_1
X_22966_ net21 VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__buf_2
XFILLER_167_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24705_ _09636_ registers\[55\]\[58\] _10569_ VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__mux2_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28473_ _11828_ registers\[28\]\[47\] _12621_ VGND VGND VPWR VPWR _12629_ sky130_fd_sc_hd__mux2_1
X_21917_ _08267_ _08579_ _08580_ _08270_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__a22o_1
X_25685_ registers\[48\]\[39\] _10386_ _11119_ VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__mux2_1
X_22897_ _09526_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27424_ registers\[36\]\[63\] _10436_ _12006_ VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24636_ _09567_ registers\[55\]\[25\] _10536_ VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__mux2_1
XFILLER_230_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21848_ registers\[0\]\[33\] registers\[1\]\[33\] registers\[2\]\[33\] registers\[3\]\[33\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__mux4_1
XFILLER_31_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_247_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27355_ _12006_ VGND VGND VPWR VPWR _12040_ sky130_fd_sc_hd__buf_4
X_24567_ _09636_ registers\[56\]\[58\] _10495_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__mux2_1
XFILLER_208_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21779_ registers\[8\]\[31\] registers\[9\]\[31\] registers\[10\]\[31\] registers\[11\]\[31\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__mux4_1
X_26306_ _10756_ registers\[43\]\[12\] _11454_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__mux2_1
X_23518_ _09605_ registers\[19\]\[43\] _09914_ VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27286_ _12003_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_211_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24498_ _09567_ registers\[56\]\[25\] _10462_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__mux2_1
X_29025_ _12919_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26237_ _11420_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23449_ _09535_ registers\[19\]\[10\] _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__mux2_1
XFILLER_99_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26168_ _11384_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25119_ net36 VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__buf_2
X_26099_ _10819_ registers\[45\]\[42\] _11345_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__mux2_1
X_18990_ registers\[20\]\[17\] registers\[21\]\[17\] registers\[22\]\[17\] registers\[23\]\[17\]
+ _05503_ _05504_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__mux4_1
XFILLER_124_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _04676_ _04713_ _04714_ _04681_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__a22o_1
X_29927_ _13425_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__clkbuf_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17872_ registers\[32\]\[51\] registers\[33\]\[51\] registers\[34\]\[51\] registers\[35\]\[51\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__mux4_1
XFILLER_152_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29858_ registers\[18\]\[32\] _13002_ _13386_ VGND VGND VPWR VPWR _13389_ sky130_fd_sc_hd__mux2_1
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19611_ _06098_ _06337_ _06338_ _06102_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a22o_1
X_28809_ _11759_ registers\[25\]\[14\] _12801_ VGND VGND VPWR VPWR _12806_ sky130_fd_sc_hd__mux2_1
X_16823_ registers\[52\]\[21\] registers\[53\]\[21\] registers\[54\]\[21\] registers\[55\]\[21\]
+ _15134_ _15135_ VGND VGND VPWR VPWR _15316_ sky130_fd_sc_hd__mux4_1
XFILLER_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_947 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29789_ _12933_ _12149_ VGND VGND VPWR VPWR _13352_ sky130_fd_sc_hd__nor2_8
XFILLER_94_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31820_ _14421_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__clkbuf_1
X_19542_ _06090_ _06270_ _06271_ _06096_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a22o_1
XFILLER_19_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16754_ registers\[12\]\[19\] registers\[13\]\[19\] registers\[14\]\[19\] registers\[15\]\[19\]
+ _15045_ _15046_ VGND VGND VPWR VPWR _15249_ sky130_fd_sc_hd__mux4_1
XFILLER_219_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_235_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19473_ registers\[48\]\[31\] registers\[49\]\[31\] registers\[50\]\[31\] registers\[51\]\[31\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__mux4_1
X_16685_ _15178_ _15181_ _14945_ VGND VGND VPWR VPWR _15182_ sky130_fd_sc_hd__o21ba_1
X_31751_ registers\[59\]\[33\] net27 _14381_ VGND VGND VPWR VPWR _14385_ sky130_fd_sc_hd__mux2_1
XFILLER_59_1157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18424_ registers\[4\]\[1\] registers\[5\]\[1\] registers\[6\]\[1\] registers\[7\]\[1\]
+ _05126_ _05128_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__mux4_1
XFILLER_181_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30702_ registers\[12\]\[48\] _13035_ _13824_ VGND VGND VPWR VPWR _13833_ sky130_fd_sc_hd__mux2_1
XFILLER_181_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34470_ clknet_leaf_464_CLK _02584_ VGND VGND VPWR VPWR registers\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31682_ registers\[59\]\[0\] net1 _14348_ VGND VGND VPWR VPWR _14349_ sky130_fd_sc_hd__mux2_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33421_ clknet_leaf_172_CLK _01535_ VGND VGND VPWR VPWR registers\[46\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_18355_ _05107_ _05110_ _05115_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__a22o_1
X_30633_ registers\[12\]\[15\] _12966_ _13791_ VGND VGND VPWR VPWR _13797_ sky130_fd_sc_hd__mux2_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ registers\[56\]\[35\] registers\[57\]\[35\] registers\[58\]\[35\] registers\[59\]\[35\]
+ _15752_ _15542_ VGND VGND VPWR VPWR _15785_ sky130_fd_sc_hd__mux4_1
X_36140_ clknet_leaf_372_CLK _04254_ VGND VGND VPWR VPWR registers\[49\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33352_ clknet_leaf_250_CLK _01466_ VGND VGND VPWR VPWR registers\[47\]\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30564_ _13760_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__clkbuf_1
X_18286_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__buf_12
XFILLER_175_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32303_ clknet_leaf_394_CLK _00417_ VGND VGND VPWR VPWR registers\[19\]\[33\] sky130_fd_sc_hd__dfxtp_1
X_17237_ registers\[36\]\[33\] registers\[37\]\[33\] registers\[38\]\[33\] registers\[39\]\[33\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15718_ sky130_fd_sc_hd__mux4_1
X_36071_ clknet_leaf_437_CLK _04185_ VGND VGND VPWR VPWR registers\[59\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_33283_ clknet_leaf_270_CLK _01397_ VGND VGND VPWR VPWR registers\[48\]\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30495_ _13724_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35022_ clknet_leaf_116_CLK _03136_ VGND VGND VPWR VPWR registers\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32234_ clknet_leaf_424_CLK _00348_ VGND VGND VPWR VPWR registers\[39\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_17168_ registers\[44\]\[31\] registers\[45\]\[31\] registers\[46\]\[31\] registers\[47\]\[31\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15651_ sky130_fd_sc_hd__mux4_2
XFILLER_156_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16119_ _14628_ _14631_ _14554_ _14556_ VGND VGND VPWR VPWR _14632_ sky130_fd_sc_hd__o211a_1
X_32165_ clknet_leaf_135_CLK _00279_ VGND VGND VPWR VPWR registers\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_963 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17099_ _15541_ _15582_ _15583_ _15547_ VGND VGND VPWR VPWR _15584_ sky130_fd_sc_hd__a22o_1
XFILLER_66_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31116_ registers\[0\]\[52\] _13044_ _14048_ VGND VGND VPWR VPWR _14051_ sky130_fd_sc_hd__mux2_1
XFILLER_192_1158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32096_ clknet_leaf_485_CLK _00009_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35924_ clknet_leaf_82_CLK _04038_ VGND VGND VPWR VPWR registers\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31047_ _14014_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19809_ _05079_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__buf_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35855_ clknet_leaf_170_CLK _03969_ VGND VGND VPWR VPWR registers\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_226_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22820_ _07325_ _09455_ _09456_ _07336_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__a22o_1
X_34806_ clknet_leaf_313_CLK _02920_ VGND VGND VPWR VPWR registers\[24\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_35786_ clknet_leaf_153_CLK _03900_ VGND VGND VPWR VPWR registers\[0\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_32998_ clknet_leaf_438_CLK _01112_ VGND VGND VPWR VPWR registers\[52\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_225_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_241_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22751_ _09109_ _09389_ _09390_ _09114_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__a22o_1
X_34737_ clknet_leaf_410_CLK _02851_ VGND VGND VPWR VPWR registers\[25\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_31949_ _14488_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21702_ _08334_ _08370_ _08371_ _08338_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__a22o_1
XFILLER_225_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25470_ registers\[4\]\[2\] _10309_ _11012_ VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__mux2_1
XFILLER_164_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22682_ registers\[12\]\[57\] registers\[13\]\[57\] registers\[14\]\[57\] registers\[15\]\[57\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__mux4_1
XFILLER_212_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34668_ clknet_leaf_410_CLK _02782_ VGND VGND VPWR VPWR registers\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_240_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24421_ _10423_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33619_ clknet_leaf_127_CLK _01733_ VGND VGND VPWR VPWR registers\[42\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_21633_ registers\[0\]\[27\] registers\[1\]\[27\] registers\[2\]\[27\] registers\[3\]\[27\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__mux4_1
XFILLER_90_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34599_ clknet_leaf_455_CLK _02713_ VGND VGND VPWR VPWR registers\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_27140_ _11847_ registers\[38\]\[56\] _11920_ VGND VGND VPWR VPWR _11927_ sky130_fd_sc_hd__mux2_1
XFILLER_139_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_240_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24352_ registers\[57\]\[34\] _10376_ _10368_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__mux2_1
XFILLER_205_1257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21564_ _07924_ _08236_ _08237_ _07927_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__a22o_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23303_ net46 VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__buf_4
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20515_ registers\[40\]\[62\] registers\[41\]\[62\] registers\[42\]\[62\] registers\[43\]\[62\]
+ _05083_ _05084_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__mux4_1
X_27071_ _11778_ registers\[38\]\[23\] _11887_ VGND VGND VPWR VPWR _11891_ sky130_fd_sc_hd__mux2_1
X_24283_ net4 VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__buf_4
X_21495_ registers\[0\]\[23\] registers\[1\]\[23\] registers\[2\]\[23\] registers\[3\]\[23\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__mux4_1
XFILLER_193_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26022_ _11307_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23234_ net22 VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20446_ registers\[24\]\[59\] registers\[25\]\[59\] registers\[26\]\[59\] registers\[27\]\[59\]
+ _07003_ _07004_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__mux4_1
XFILLER_119_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23165_ registers\[9\]\[2\] _09662_ _09709_ VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__mux2_1
XFILLER_162_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20377_ _06784_ _07081_ _07082_ _06788_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__a22o_1
XTAP_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22116_ _08741_ _08750_ _08760_ _08774_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__or4_4
XTAP_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27973_ _12366_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__clkbuf_1
X_23096_ net34 VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__buf_4
XANTENNA_1209 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29712_ registers\[1\]\[27\] _12991_ _13304_ VGND VGND VPWR VPWR _13312_ sky130_fd_sc_hd__mux2_1
XTAP_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26924_ _11798_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22047_ registers\[36\]\[39\] registers\[37\]\[39\] registers\[38\]\[39\] registers\[39\]\[39\]
+ _08635_ _08636_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__mux4_1
XFILLER_248_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1091 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29643_ _13275_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__clkbuf_1
XTAP_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26855_ _11750_ registers\[3\]\[10\] _11751_ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__mux2_1
XTAP_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_25806_ _10796_ registers\[47\]\[31\] _11192_ VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__mux2_1
X_26786_ registers\[40\]\[47\] _10403_ _11702_ VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__mux2_1
X_29574_ _13239_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23998_ _09538_ registers\[5\]\[11\] _10172_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__mux2_1
X_25737_ net87 _09650_ net88 VGND VGND VPWR VPWR _11156_ sky130_fd_sc_hd__and3b_1
X_28525_ _12656_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22949_ _09561_ registers\[62\]\[22\] _09557_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__mux2_1
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16470_ registers\[52\]\[11\] registers\[53\]\[11\] registers\[54\]\[11\] registers\[55\]\[11\]
+ _14791_ _14792_ VGND VGND VPWR VPWR _14973_ sky130_fd_sc_hd__mux4_1
X_25668_ _11120_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
X_28456_ _11811_ registers\[28\]\[39\] _12610_ VGND VGND VPWR VPWR _12620_ sky130_fd_sc_hd__mux2_1
XFILLER_243_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27407_ _12067_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24619_ _09550_ registers\[55\]\[17\] _10525_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__mux2_1
X_28387_ _11742_ registers\[28\]\[6\] _12577_ VGND VGND VPWR VPWR _12584_ sky130_fd_sc_hd__mux2_1
X_25599_ _10512_ VGND VGND VPWR VPWR _11082_ sky130_fd_sc_hd__inv_2
XFILLER_169_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18140_ registers\[0\]\[59\] registers\[1\]\[59\] registers\[2\]\[59\] registers\[3\]\[59\]
+ _04623_ _04624_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__mux4_1
XFILLER_157_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27338_ _12031_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18071_ _04837_ _04840_ _04611_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__o21ba_2
X_27269_ _11841_ registers\[37\]\[53\] _11991_ VGND VGND VPWR VPWR _11995_ sky130_fd_sc_hd__mux2_1
XFILLER_157_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17022_ registers\[36\]\[27\] registers\[37\]\[27\] registers\[38\]\[27\] registers\[39\]\[27\]
+ _15507_ _15508_ VGND VGND VPWR VPWR _15509_ sky130_fd_sc_hd__mux4_1
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29008_ _12910_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30280_ registers\[15\]\[40\] _13018_ _13610_ VGND VGND VPWR VPWR _13611_ sky130_fd_sc_hd__mux2_1
XFILLER_236_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18973_ registers\[48\]\[17\] registers\[49\]\[17\] registers\[50\]\[17\] registers\[51\]\[17\]
+ _05407_ _05408_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__mux4_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1710 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1721 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ registers\[12\]\[52\] registers\[13\]\[52\] registers\[14\]\[52\] registers\[15\]\[52\]
+ _04387_ _04388_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux4_1
XANTENNA_1732 _00178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1743 _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33970_ clknet_leaf_356_CLK _02084_ VGND VGND VPWR VPWR registers\[37\]\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1754 _07295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1765 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32921_ clknet_leaf_62_CLK _01035_ VGND VGND VPWR VPWR registers\[53\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1776 _11864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ _14490_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1787 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35640_ clknet_leaf_317_CLK _03754_ VGND VGND VPWR VPWR registers\[11\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_16806_ _14610_ VGND VGND VPWR VPWR _15300_ sky130_fd_sc_hd__clkbuf_4
X_32852_ clknet_leaf_64_CLK _00966_ VGND VGND VPWR VPWR registers\[54\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_17786_ registers\[16\]\[48\] registers\[17\]\[48\] registers\[18\]\[48\] registers\[19\]\[48\]
+ _04493_ _04494_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__mux4_1
X_31803_ registers\[59\]\[58\] net54 _14403_ VGND VGND VPWR VPWR _14412_ sky130_fd_sc_hd__mux2_1
X_19525_ _05125_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__buf_6
XFILLER_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35571_ clknet_leaf_354_CLK _03685_ VGND VGND VPWR VPWR registers\[12\]\[37\] sky130_fd_sc_hd__dfxtp_1
X_16737_ _14520_ VGND VGND VPWR VPWR _15232_ sky130_fd_sc_hd__buf_4
X_32783_ clknet_leaf_173_CLK _00897_ VGND VGND VPWR VPWR registers\[55\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34522_ clknet_leaf_3_CLK _02636_ VGND VGND VPWR VPWR registers\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19456_ _05079_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__buf_4
X_31734_ registers\[59\]\[25\] net18 _14370_ VGND VGND VPWR VPWR _14376_ sky130_fd_sc_hd__mux2_1
XFILLER_201_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16668_ _14573_ VGND VGND VPWR VPWR _15165_ sky130_fd_sc_hd__buf_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_228_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18407_ registers\[44\]\[1\] registers\[45\]\[1\] registers\[46\]\[1\] registers\[47\]\[1\]
+ _05061_ _05062_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__mux4_1
XFILLER_37_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34453_ clknet_leaf_80_CLK _02567_ VGND VGND VPWR VPWR registers\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_222_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31665_ _14339_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__clkbuf_1
X_19387_ _06121_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16599_ _15094_ _15097_ _14926_ VGND VGND VPWR VPWR _15098_ sky130_fd_sc_hd__o21ba_1
X_33404_ clknet_leaf_278_CLK _01518_ VGND VGND VPWR VPWR registers\[46\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_18338_ _05089_ _05094_ _05099_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a22o_1
X_30616_ registers\[12\]\[7\] _12949_ _13780_ VGND VGND VPWR VPWR _13788_ sky130_fd_sc_hd__mux2_1
XFILLER_241_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34384_ clknet_leaf_100_CLK _02498_ VGND VGND VPWR VPWR registers\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_31596_ _14303_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__clkbuf_1
X_36123_ clknet_leaf_36_CLK _04237_ VGND VGND VPWR VPWR registers\[49\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_33335_ clknet_leaf_342_CLK _01449_ VGND VGND VPWR VPWR registers\[47\]\[41\] sky130_fd_sc_hd__dfxtp_1
X_18269_ registers\[28\]\[63\] registers\[29\]\[63\] registers\[30\]\[63\] registers\[31\]\[63\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__mux4_1
X_30547_ _13751_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20300_ registers\[20\]\[54\] registers\[21\]\[54\] registers\[22\]\[54\] registers\[23\]\[54\]
+ _06875_ _06876_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__mux4_1
XFILLER_159_1318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36054_ clknet_leaf_67_CLK _04168_ VGND VGND VPWR VPWR registers\[59\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21280_ registers\[0\]\[17\] registers\[1\]\[17\] registers\[2\]\[17\] registers\[3\]\[17\]
+ _07723_ _07724_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__mux4_1
X_33266_ clknet_leaf_364_CLK _01380_ VGND VGND VPWR VPWR registers\[48\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_30478_ _13715_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35005_ clknet_leaf_186_CLK _03119_ VGND VGND VPWR VPWR registers\[21\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20231_ _05125_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__buf_6
X_32217_ clknet_leaf_295_CLK _00331_ VGND VGND VPWR VPWR registers\[9\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33197_ clknet_leaf_390_CLK _01311_ VGND VGND VPWR VPWR registers\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_239_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20162_ _05079_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__buf_4
XFILLER_171_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32148_ clknet_leaf_119_CLK _00262_ VGND VGND VPWR VPWR registers\[39\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24970_ _10718_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__clkbuf_1
X_20093_ _06807_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
X_32079_ clknet_leaf_491_CLK _00011_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dfxtp_1
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23921_ _10132_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
X_35907_ clknet_leaf_233_CLK _04021_ VGND VGND VPWR VPWR registers\[7\]\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_893 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26640_ _10819_ registers\[41\]\[42\] _11630_ VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__mux2_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35838_ clknet_leaf_295_CLK _03952_ VGND VGND VPWR VPWR registers\[8\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_23852_ _10096_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__clkbuf_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22803_ registers\[4\]\[61\] registers\[5\]\[61\] registers\[6\]\[61\] registers\[7\]\[61\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__mux4_1
XANTENNA_607 _05104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26571_ _11596_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__clkbuf_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35769_ clknet_leaf_316_CLK _03883_ VGND VGND VPWR VPWR registers\[0\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_23783_ _10059_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__clkbuf_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_618 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20995_ registers\[52\]\[9\] registers\[53\]\[9\] registers\[54\]\[9\] registers\[55\]\[9\]
+ _07576_ _07577_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__mux4_1
XANTENNA_629 _05127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28310_ _12543_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__clkbuf_1
X_25522_ registers\[4\]\[27\] _10361_ _11034_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22734_ _07372_ _09372_ _09373_ _07382_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__a22o_1
X_29290_ _09697_ registers\[22\]\[19\] _13080_ VGND VGND VPWR VPWR _13090_ sky130_fd_sc_hd__mux2_1
XFILLER_214_967 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_1319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28241_ _12507_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25453_ _11003_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1057 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22665_ registers\[40\]\[57\] registers\[41\]\[57\] registers\[42\]\[57\] registers\[43\]\[57\]
+ _09149_ _09150_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__mux4_1
XFILLER_241_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24404_ net47 VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__buf_4
XFILLER_240_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28172_ _11797_ registers\[30\]\[32\] _12468_ VGND VGND VPWR VPWR _12471_ sky130_fd_sc_hd__mux2_1
X_21616_ registers\[40\]\[27\] registers\[41\]\[27\] registers\[42\]\[27\] registers\[43\]\[27\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__mux4_1
XFILLER_107_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25384_ _10967_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__clkbuf_1
X_22596_ registers\[24\]\[54\] registers\[25\]\[54\] registers\[26\]\[54\] registers\[27\]\[54\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__mux4_1
XFILLER_187_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27123_ _11830_ registers\[38\]\[48\] _11909_ VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__mux2_1
XFILLER_16_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24335_ net22 VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__buf_4
X_21547_ registers\[32\]\[25\] registers\[33\]\[25\] registers\[34\]\[25\] registers\[35\]\[25\]
+ _08016_ _08017_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__mux4_1
XFILLER_14_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27054_ _11761_ registers\[38\]\[15\] _11876_ VGND VGND VPWR VPWR _11882_ sky130_fd_sc_hd__mux2_1
XFILLER_166_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24266_ _10318_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21478_ _08131_ _08138_ _08145_ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__or4_4
XFILLER_107_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26005_ _10860_ registers\[46\]\[62\] _11229_ VGND VGND VPWR VPWR _11298_ sky130_fd_sc_hd__mux2_1
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23217_ net17 VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20429_ registers\[36\]\[59\] registers\[37\]\[59\] registers\[38\]\[59\] registers\[39\]\[59\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__mux4_1
XFILLER_84_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24197_ _09601_ registers\[58\]\[41\] _10277_ VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__mux2_1
XFILLER_101_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23148_ net13 VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__clkbuf_4
XTAP_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1006 _11843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1017 _12363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1028 _12934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23079_ net86 VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__clkbuf_4
X_27956_ registers\[32\]\[58\] _10426_ _12348_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__mux2_1
XTAP_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1039 _13139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26907_ _11786_ registers\[3\]\[27\] _11772_ VGND VGND VPWR VPWR _11787_ sky130_fd_sc_hd__mux2_1
XFILLER_248_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27887_ registers\[32\]\[25\] _10357_ _12315_ VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__mux2_1
XTAP_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29626_ registers\[20\]\[50\] _13039_ _13266_ VGND VGND VPWR VPWR _13267_ sky130_fd_sc_hd__mux2_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _04419_ _04422_ _15974_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o21ba_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26838_ net56 VGND VGND VPWR VPWR _11740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29557_ _13230_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17571_ registers\[12\]\[42\] registers\[13\]\[42\] registers\[14\]\[42\] registers\[15\]\[42\]
+ _15731_ _15732_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__mux4_1
X_26769_ registers\[40\]\[39\] _10386_ _11691_ VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__mux2_1
XFILLER_95_1132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19310_ registers\[28\]\[26\] registers\[29\]\[26\] registers\[30\]\[26\] registers\[31\]\[26\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__mux4_1
X_28508_ _09868_ _10014_ VGND VGND VPWR VPWR _12647_ sky130_fd_sc_hd__nand2_8
X_16522_ registers\[20\]\[12\] registers\[21\]\[12\] registers\[22\]\[12\] registers\[23\]\[12\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _15024_ sky130_fd_sc_hd__mux4_1
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29488_ _09795_ registers\[21\]\[49\] _13184_ VGND VGND VPWR VPWR _13194_ sky130_fd_sc_hd__mux2_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19241_ registers\[20\]\[24\] registers\[21\]\[24\] registers\[22\]\[24\] registers\[23\]\[24\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__mux4_1
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_1198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28439_ _12611_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__clkbuf_1
X_16453_ _14610_ VGND VGND VPWR VPWR _14957_ sky130_fd_sc_hd__clkbuf_4
XFILLER_231_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_220_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_223_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_959 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16384_ _14520_ VGND VGND VPWR VPWR _14889_ sky130_fd_sc_hd__clkbuf_8
X_31450_ _14226_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__clkbuf_1
X_19172_ _05141_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__buf_4
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18123_ _04870_ _04877_ _04884_ _04891_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__or4_4
XFILLER_185_852 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30401_ _09760_ registers\[14\]\[33\] _13671_ VGND VGND VPWR VPWR _13675_ sky130_fd_sc_hd__mux2_1
X_31381_ _14134_ VGND VGND VPWR VPWR _14190_ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_1417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_200_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33120_ clknet_leaf_42_CLK _01234_ VGND VGND VPWR VPWR registers\[50\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_18054_ _14511_ _04823_ _04824_ _14517_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a22o_1
X_30332_ _09648_ registers\[14\]\[0\] _13638_ VGND VGND VPWR VPWR _13639_ sky130_fd_sc_hd__mux2_1
XFILLER_144_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17005_ registers\[24\]\[26\] registers\[25\]\[26\] registers\[26\]\[26\] registers\[27\]\[26\]
+ _15425_ _15426_ VGND VGND VPWR VPWR _15493_ sky130_fd_sc_hd__mux4_1
X_33051_ clknet_leaf_35_CLK _01165_ VGND VGND VPWR VPWR registers\[51\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_30263_ registers\[15\]\[32\] _13002_ _13599_ VGND VGND VPWR VPWR _13602_ sky130_fd_sc_hd__mux2_1
XFILLER_119_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32002_ clknet_leaf_27_CLK _00175_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
X_30194_ _09656_ _09705_ VGND VGND VPWR VPWR _13565_ sky130_fd_sc_hd__nor2_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18956_ _05496_ _05699_ _05702_ _05499_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__a22o_1
XANTENNA_1540 _09793_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1551 _11300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17907_ _04676_ _04679_ _04680_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a22o_1
XFILLER_234_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1562 _11748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33953_ clknet_leaf_41_CLK _02067_ VGND VGND VPWR VPWR registers\[37\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1573 _13068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18887_ registers\[28\]\[14\] registers\[29\]\[14\] registers\[30\]\[14\] registers\[31\]\[14\]
+ _05570_ _05571_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__mux4_1
XFILLER_39_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_230_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1584 _14489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1595 _14548_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32904_ clknet_leaf_178_CLK _01018_ VGND VGND VPWR VPWR registers\[54\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_17838_ _04540_ _04613_ _04614_ _04546_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__a22o_1
XFILLER_27_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33884_ clknet_leaf_23_CLK _01998_ VGND VGND VPWR VPWR registers\[38\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35623_ clknet_leaf_460_CLK _03737_ VGND VGND VPWR VPWR registers\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_208_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32835_ clknet_leaf_293_CLK _00949_ VGND VGND VPWR VPWR registers\[55\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_17769_ _14509_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__buf_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19508_ registers\[56\]\[32\] registers\[57\]\[32\] registers\[58\]\[32\] registers\[59\]\[32\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__mux4_1
XFILLER_78_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35554_ clknet_leaf_467_CLK _03668_ VGND VGND VPWR VPWR registers\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20780_ _07472_ _07475_ _07310_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__o21ba_1
X_32766_ clknet_leaf_291_CLK _00880_ VGND VGND VPWR VPWR registers\[56\]\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34505_ clknet_leaf_217_CLK _02619_ VGND VGND VPWR VPWR registers\[2\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_19439_ registers\[8\]\[30\] registers\[9\]\[30\] registers\[10\]\[30\] registers\[11\]\[30\]
+ _05998_ _05999_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__mux4_1
X_31717_ registers\[59\]\[17\] net9 _14359_ VGND VGND VPWR VPWR _14367_ sky130_fd_sc_hd__mux2_1
X_35485_ clknet_leaf_482_CLK _03599_ VGND VGND VPWR VPWR registers\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_223_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32697_ clknet_leaf_333_CLK _00811_ VGND VGND VPWR VPWR registers\[57\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_245_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22450_ registers\[12\]\[50\] registers\[13\]\[50\] registers\[14\]\[50\] registers\[15\]\[50\]
+ _08859_ _08860_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__mux4_1
X_34436_ clknet_leaf_206_CLK _02550_ VGND VGND VPWR VPWR registers\[30\]\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31648_ _14330_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_241_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21401_ _07385_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__clkbuf_4
X_22381_ _07363_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__buf_4
X_34367_ clknet_leaf_188_CLK _02481_ VGND VGND VPWR VPWR registers\[31\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31579_ _14294_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_822 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36106_ clknet_leaf_176_CLK _04220_ VGND VGND VPWR VPWR registers\[59\]\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24120_ _10238_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__clkbuf_1
X_33318_ clknet_leaf_61_CLK _01432_ VGND VGND VPWR VPWR registers\[47\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_21332_ _08009_ _08012_ _07744_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__o21ba_1
X_34298_ clknet_leaf_280_CLK _02412_ VGND VGND VPWR VPWR registers\[32\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36037_ clknet_leaf_199_CLK _04151_ VGND VGND VPWR VPWR registers\[63\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24051_ _10201_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33249_ clknet_leaf_42_CLK _01363_ VGND VGND VPWR VPWR registers\[48\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_21263_ registers\[40\]\[17\] registers\[41\]\[17\] registers\[42\]\[17\] registers\[43\]\[17\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__mux4_1
XFILLER_190_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23002_ _09597_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_20214_ registers\[56\]\[52\] registers\[57\]\[52\] registers\[58\]\[52\] registers\[59\]\[52\]
+ _06644_ _06777_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__mux4_1
XFILLER_172_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap283 _10304_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21194_ registers\[32\]\[15\] registers\[33\]\[15\] registers\[34\]\[15\] registers\[35\]\[15\]
+ _07673_ _07674_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27810_ _12280_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__clkbuf_1
X_20145_ registers\[8\]\[50\] registers\[9\]\[50\] registers\[10\]\[50\] registers\[11\]\[50\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__mux4_1
X_28790_ _11740_ registers\[25\]\[5\] _12790_ VGND VGND VPWR VPWR _12796_ sky130_fd_sc_hd__mux2_1
XFILLER_246_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24953_ _10709_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__clkbuf_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27741_ _12221_ VGND VGND VPWR VPWR _12244_ sky130_fd_sc_hd__buf_4
XFILLER_170_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20076_ registers\[8\]\[48\] registers\[9\]\[48\] registers\[10\]\[48\] registers\[11\]\[48\]
+ _06684_ _06685_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__mux4_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23904_ _09580_ registers\[60\]\[31\] _10122_ VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__mux2_1
XFILLER_245_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27672_ registers\[34\]\[51\] _10412_ _12206_ VGND VGND VPWR VPWR _12208_ sky130_fd_sc_hd__mux2_1
X_24884_ _10673_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__clkbuf_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_246_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29411_ _09683_ registers\[21\]\[12\] _13151_ VGND VGND VPWR VPWR _13154_ sky130_fd_sc_hd__mux2_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23835_ _10086_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
X_26623_ _10802_ registers\[41\]\[34\] _11619_ VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__mux2_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_404 _00096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_415 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_426 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26554_ _10733_ registers\[41\]\[1\] _11586_ VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__mux2_1
XANTENNA_437 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_29342_ _13117_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23766_ _09577_ registers\[29\]\[30\] _10050_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__mux2_1
XANTENNA_448 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20978_ _07386_ _07667_ _07668_ _07396_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__a22o_1
XANTENNA_459 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22717_ registers\[16\]\[58\] registers\[17\]\[58\] registers\[18\]\[58\] registers\[19\]\[58\]
+ _07387_ _07389_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__mux4_1
X_25505_ registers\[4\]\[19\] _10344_ _11023_ VGND VGND VPWR VPWR _11033_ sky130_fd_sc_hd__mux2_1
XFILLER_144_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29273_ _13081_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__clkbuf_1
X_26485_ _10800_ registers\[42\]\[33\] _11547_ VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__mux2_1
X_23697_ _10012_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28224_ _11849_ registers\[30\]\[57\] _12490_ VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__mux2_1
X_25436_ _10840_ registers\[50\]\[52\] _10992_ VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__mux2_1
XFILLER_158_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22648_ _09287_ _09290_ _09091_ _09092_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__o211a_1
XFILLER_224_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_194_CLK clknet_6_49__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_194_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_28155_ _11780_ registers\[30\]\[24\] _12457_ VGND VGND VPWR VPWR _12462_ sky130_fd_sc_hd__mux2_1
X_25367_ _10958_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_210_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22579_ registers\[56\]\[54\] registers\[57\]\[54\] registers\[58\]\[54\] registers\[59\]\[54\]
+ _09223_ _09013_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__mux4_1
X_27106_ _11864_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__buf_4
X_24318_ registers\[57\]\[23\] _10353_ _10347_ VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__mux2_1
X_28086_ _12425_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__clkbuf_1
X_25298_ _10838_ registers\[51\]\[51\] _10920_ VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__mux2_1
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27037_ _11744_ registers\[38\]\[7\] _11865_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__mux2_1
X_24249_ net12 VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_1404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_218_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18810_ registers\[0\]\[12\] registers\[1\]\[12\] registers\[2\]\[12\] registers\[3\]\[12\]
+ _05487_ _05488_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__mux4_1
XTAP_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19790_ _05104_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28988_ registers\[24\]\[35\] _10378_ _12894_ VGND VGND VPWR VPWR _12900_ sky130_fd_sc_hd__mux2_1
XTAP_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput95 net95 VGND VGND VPWR VPWR D1[14] sky130_fd_sc_hd__buf_2
XTAP_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18741_ _05133_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__buf_2
X_27939_ _12292_ VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__buf_4
XTAP_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18672_ _05421_ _05426_ _05134_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__o21ba_1
X_30950_ _13963_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__clkbuf_1
XTAP_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _04340_ _04404_ _04405_ _04343_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__a22o_1
X_29609_ registers\[20\]\[42\] _13023_ _13255_ VGND VGND VPWR VPWR _13258_ sky130_fd_sc_hd__mux2_1
XFILLER_224_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_30881_ _13927_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__clkbuf_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_236_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_229_1330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_32620_ clknet_leaf_372_CLK _00734_ VGND VGND VPWR VPWR registers\[58\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _04333_ _04336_ _04337_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a22o_1
XFILLER_204_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_232_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_960 _10836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_220_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_971 _11085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16505_ registers\[60\]\[12\] registers\[61\]\[12\] registers\[62\]\[12\] registers\[63\]\[12\]
+ _14727_ _14864_ VGND VGND VPWR VPWR _15007_ sky130_fd_sc_hd__mux4_1
X_32551_ clknet_leaf_457_CLK _00665_ VGND VGND VPWR VPWR registers\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_982 _11300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17485_ _15884_ _15957_ _15958_ _15890_ VGND VGND VPWR VPWR _15959_ sky130_fd_sc_hd__a22o_1
XANTENNA_993 _11755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_204_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31502_ _09782_ registers\[6\]\[43\] _14250_ VGND VGND VPWR VPWR _14254_ sky130_fd_sc_hd__mux2_1
X_19224_ registers\[60\]\[24\] registers\[61\]\[24\] registers\[62\]\[24\] registers\[63\]\[24\]
+ _05962_ _05756_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__mux4_1
X_35270_ clknet_leaf_154_CLK _03384_ VGND VGND VPWR VPWR registers\[17\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_177_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16436_ registers\[0\]\[10\] registers\[1\]\[10\] registers\[2\]\[10\] registers\[3\]\[10\]
+ _14938_ _14939_ VGND VGND VPWR VPWR _14940_ sky130_fd_sc_hd__mux4_1
X_32482_ clknet_leaf_444_CLK _00596_ VGND VGND VPWR VPWR registers\[60\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34221_ clknet_leaf_321_CLK _02335_ VGND VGND VPWR VPWR registers\[33\]\[31\] sky130_fd_sc_hd__dfxtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31433_ _09678_ registers\[6\]\[10\] _14217_ VGND VGND VPWR VPWR _14218_ sky130_fd_sc_hd__mux2_1
X_19155_ registers\[56\]\[22\] registers\[57\]\[22\] registers\[58\]\[22\] registers\[59\]\[22\]
+ _05615_ _05748_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__mux4_1
X_16367_ registers\[12\]\[8\] registers\[13\]\[8\] registers\[14\]\[8\] registers\[15\]\[8\]
+ _14702_ _14703_ VGND VGND VPWR VPWR _14873_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_185_CLK clknet_6_48__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_185_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18106_ registers\[52\]\[58\] registers\[53\]\[58\] registers\[54\]\[58\] registers\[55\]\[58\]
+ _14494_ _14497_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__mux4_1
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34152_ clknet_leaf_431_CLK _02266_ VGND VGND VPWR VPWR registers\[34\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16298_ _14800_ _14805_ _14585_ VGND VGND VPWR VPWR _14806_ sky130_fd_sc_hd__o21ba_1
XFILLER_121_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19086_ registers\[8\]\[20\] registers\[9\]\[20\] registers\[10\]\[20\] registers\[11\]\[20\]
+ _05655_ _05656_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__mux4_1
X_31364_ _14181_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33103_ clknet_leaf_75_CLK _01217_ VGND VGND VPWR VPWR registers\[50\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_18037_ _04676_ _04806_ _04807_ _04681_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__a22o_1
X_30315_ registers\[15\]\[57\] _13054_ _13621_ VGND VGND VPWR VPWR _13629_ sky130_fd_sc_hd__mux2_1
XFILLER_219_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_6_33__f_CLK clknet_5_16_0_CLK VGND VGND VPWR VPWR clknet_6_33__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_34083_ clknet_leaf_47_CLK _02197_ VGND VGND VPWR VPWR registers\[35\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31295_ registers\[7\]\[9\] net64 _14135_ VGND VGND VPWR VPWR _14145_ sky130_fd_sc_hd__mux2_1
XFILLER_160_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_33034_ clknet_leaf_162_CLK _01148_ VGND VGND VPWR VPWR registers\[52\]\[60\] sky130_fd_sc_hd__dfxtp_1
X_30246_ registers\[15\]\[24\] _12985_ _13588_ VGND VGND VPWR VPWR _13593_ sky130_fd_sc_hd__mux2_1
XFILLER_99_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30177_ _13556_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__clkbuf_1
X_19988_ registers\[36\]\[46\] registers\[37\]\[46\] registers\[38\]\[46\] registers\[39\]\[46\]
+ _06399_ _06400_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux4_1
XFILLER_132_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18939_ _05412_ _05682_ _05685_ _05416_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__a22o_1
XFILLER_189_1108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34985_ clknet_leaf_453_CLK _03099_ VGND VGND VPWR VPWR registers\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1370 _00170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1381 _00171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_223_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33936_ clknet_leaf_121_CLK _02050_ VGND VGND VPWR VPWR registers\[37\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1392 _00172_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21950_ _07352_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__buf_4
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20901_ _07379_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__buf_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33867_ clknet_leaf_151_CLK _01981_ VGND VGND VPWR VPWR registers\[3\]\[61\] sky130_fd_sc_hd__dfxtp_1
X_21881_ registers\[8\]\[34\] registers\[9\]\[34\] registers\[10\]\[34\] registers\[11\]\[34\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__mux4_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35606_ clknet_leaf_86_CLK _03720_ VGND VGND VPWR VPWR registers\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23620_ _09972_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
X_20832_ registers\[16\]\[4\] registers\[17\]\[4\] registers\[18\]\[4\] registers\[19\]\[4\]
+ _07378_ _07380_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__mux4_1
X_32818_ clknet_leaf_355_CLK _00932_ VGND VGND VPWR VPWR registers\[55\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_33798_ clknet_leaf_248_CLK _01912_ VGND VGND VPWR VPWR registers\[40\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23551_ _09638_ registers\[19\]\[59\] _09925_ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__mux2_1
X_35537_ clknet_leaf_107_CLK _03651_ VGND VGND VPWR VPWR registers\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_211_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20763_ registers\[24\]\[2\] registers\[25\]\[2\] registers\[26\]\[2\] registers\[27\]\[2\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__mux4_1
XFILLER_23_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32749_ clknet_leaf_373_CLK _00863_ VGND VGND VPWR VPWR registers\[56\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22502_ _07278_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__buf_8
X_26270_ _11437_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
X_35468_ clknet_leaf_150_CLK _03582_ VGND VGND VPWR VPWR registers\[14\]\[62\] sky130_fd_sc_hd__dfxtp_1
X_23482_ _09569_ registers\[19\]\[26\] _09892_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__mux2_1
XFILLER_211_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20694_ _07392_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__buf_4
XFILLER_149_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25221_ _10881_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkbuf_1
X_22433_ _08812_ _09080_ _09081_ _08815_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__a22o_1
XFILLER_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34419_ clknet_leaf_413_CLK _02533_ VGND VGND VPWR VPWR registers\[30\]\[37\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_176_CLK clknet_6_27__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_176_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_148_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_35399_ clknet_leaf_215_CLK _03513_ VGND VGND VPWR VPWR registers\[15\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25152_ _10839_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22364_ _07326_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__buf_4
XFILLER_108_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24103_ _10228_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21315_ _07991_ _07993_ _07994_ _07995_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__a22o_1
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29960_ _13442_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__clkbuf_1
X_25083_ _10792_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
X_22295_ _07331_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__buf_4
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28911_ _11861_ registers\[25\]\[63\] _12789_ VGND VGND VPWR VPWR _12859_ sky130_fd_sc_hd__mux2_1
X_24034_ _10192_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__clkbuf_1
X_21246_ _07295_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__clkbuf_4
X_29891_ registers\[18\]\[48\] _13035_ _13397_ VGND VGND VPWR VPWR _13406_ sky130_fd_sc_hd__mux2_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_1164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_215_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28842_ _12789_ VGND VGND VPWR VPWR _12823_ sky130_fd_sc_hd__buf_4
XFILLER_89_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21177_ _07581_ _07860_ _07861_ _07584_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__a22o_1
XFILLER_120_925 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20128_ _06569_ _06839_ _06840_ _06574_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__a22o_1
X_28773_ _12786_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_213_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25985_ _10840_ registers\[46\]\[52\] _11285_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__mux2_1
XFILLER_86_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_213_1153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27724_ _12235_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_100_CLK clknet_6_17__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_100_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20059_ _06576_ _06772_ _06773_ _06579_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__a22o_1
X_24936_ _10700_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_248_1205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27655_ registers\[34\]\[43\] _10395_ _12195_ VGND VGND VPWR VPWR _12199_ sky130_fd_sc_hd__mux2_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24867_ _10664_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_201 _00053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_212 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_223 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26606_ _10785_ registers\[41\]\[26\] _11608_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__mux2_1
XFILLER_22_1192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23818_ _09630_ registers\[29\]\[55\] _10072_ VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__mux2_1
XANTENNA_234 _00056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27586_ registers\[34\]\[10\] _10325_ _12162_ VGND VGND VPWR VPWR _12163_ sky130_fd_sc_hd__mux2_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24798_ _09592_ registers\[54\]\[37\] _10620_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__mux2_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _00057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29325_ _13108_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__clkbuf_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26537_ _10852_ registers\[42\]\[58\] _11569_ VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__mux2_1
XANTENNA_278 _00058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23749_ _09561_ registers\[29\]\[22\] _10039_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__mux2_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 _00059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29256_ _13072_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17270_ _15684_ _15748_ _15749_ _15687_ VGND VGND VPWR VPWR _15750_ sky130_fd_sc_hd__a22o_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26468_ _10783_ registers\[42\]\[25\] _11536_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__mux2_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16221_ _14726_ _14730_ _14554_ _14556_ VGND VGND VPWR VPWR _14731_ sky130_fd_sc_hd__o211a_1
X_28207_ _11832_ registers\[30\]\[49\] _12479_ VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_167_CLK clknet_6_28__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_167_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_25419_ _10823_ registers\[50\]\[44\] _10981_ VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__mux2_1
X_26399_ _11505_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__clkbuf_1
X_29187_ _13026_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_201_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16152_ registers\[60\]\[2\] registers\[61\]\[2\] registers\[62\]\[2\] registers\[63\]\[2\]
+ _14542_ _14544_ VGND VGND VPWR VPWR _14664_ sky130_fd_sc_hd__mux4_1
XFILLER_31_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28138_ _11763_ registers\[30\]\[16\] _12446_ VGND VGND VPWR VPWR _12453_ sky130_fd_sc_hd__mux2_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16083_ _14499_ VGND VGND VPWR VPWR _14597_ sky130_fd_sc_hd__clkbuf_16
XFILLER_181_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28069_ _12416_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19911_ _06525_ _06629_ _06630_ _06528_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__a22o_1
X_30100_ registers\[16\]\[19\] _12974_ _13506_ VGND VGND VPWR VPWR _13516_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31080_ registers\[0\]\[35\] _13008_ _14026_ VGND VGND VPWR VPWR _14032_ sky130_fd_sc_hd__mux2_1
XFILLER_177_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_869 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30031_ registers\[17\]\[50\] _13039_ _13479_ VGND VGND VPWR VPWR _13480_ sky130_fd_sc_hd__mux2_1
XFILLER_155_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_218_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19842_ registers\[28\]\[41\] registers\[29\]\[41\] registers\[30\]\[41\] registers\[31\]\[41\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__mux4_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19773_ registers\[40\]\[40\] registers\[41\]\[40\] registers\[42\]\[40\] registers\[43\]\[40\]
+ _06227_ _06228_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__mux4_1
X_16985_ registers\[56\]\[26\] registers\[57\]\[26\] registers\[58\]\[26\] registers\[59\]\[26\]
+ _15409_ _15199_ VGND VGND VPWR VPWR _15473_ sky130_fd_sc_hd__mux4_1
XFILLER_7_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18724_ registers\[56\]\[10\] registers\[57\]\[10\] registers\[58\]\[10\] registers\[59\]\[10\]
+ _05272_ _05405_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__mux4_1
XFILLER_114_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34770_ clknet_leaf_80_CLK _02884_ VGND VGND VPWR VPWR registers\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31982_ clknet_leaf_21_CLK _00153_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_92_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33721_ clknet_leaf_338_CLK _01835_ VGND VGND VPWR VPWR registers\[41\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_18655_ _05049_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__clkbuf_4
X_30933_ _13954_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17606_ registers\[4\]\[43\] registers\[5\]\[43\] registers\[6\]\[43\] registers\[7\]\[43\]
+ _15903_ _15904_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__mux4_1
XFILLER_188_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33652_ clknet_leaf_344_CLK _01766_ VGND VGND VPWR VPWR registers\[42\]\[38\] sky130_fd_sc_hd__dfxtp_1
X_30864_ _09821_ registers\[11\]\[61\] _13850_ VGND VGND VPWR VPWR _13918_ sky130_fd_sc_hd__mux2_1
XFILLER_224_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18586_ _05089_ _05339_ _05342_ _05100_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__a22o_1
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_224_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32603_ clknet_leaf_36_CLK _00717_ VGND VGND VPWR VPWR registers\[58\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_903 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17537_ _15830_ _04321_ _04322_ _15833_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a22o_1
XFILLER_205_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33583_ clknet_leaf_360_CLK _01697_ VGND VGND VPWR VPWR registers\[43\]\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_229_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30795_ _09749_ registers\[11\]\[28\] _13873_ VGND VGND VPWR VPWR _13882_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_790 _08872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35322_ clknet_leaf_185_CLK _03436_ VGND VGND VPWR VPWR registers\[16\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32534_ clknet_leaf_68_CLK _00648_ VGND VGND VPWR VPWR registers\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17468_ registers\[20\]\[39\] registers\[21\]\[39\] registers\[22\]\[39\] registers\[23\]\[39\]
+ _15640_ _15641_ VGND VGND VPWR VPWR _15943_ sky130_fd_sc_hd__mux4_1
XFILLER_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_19207_ registers\[20\]\[23\] registers\[21\]\[23\] registers\[22\]\[23\] registers\[23\]\[23\]
+ _05846_ _05847_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__mux4_1
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16419_ registers\[44\]\[10\] registers\[45\]\[10\] registers\[46\]\[10\] registers\[47\]\[10\]
+ _14921_ _14922_ VGND VGND VPWR VPWR _14923_ sky130_fd_sc_hd__mux4_1
X_35253_ clknet_leaf_417_CLK _03367_ VGND VGND VPWR VPWR registers\[17\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_242_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_158_CLK clknet_6_31__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_158_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_32465_ clknet_leaf_179_CLK _00579_ VGND VGND VPWR VPWR registers\[60\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_220_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17399_ _15854_ _15861_ _15868_ _15875_ VGND VGND VPWR VPWR _15876_ sky130_fd_sc_hd__or4_4
XFILLER_160_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34204_ clknet_leaf_23_CLK _02318_ VGND VGND VPWR VPWR registers\[33\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_31416_ _09662_ registers\[6\]\[2\] _14206_ VGND VGND VPWR VPWR _14209_ sky130_fd_sc_hd__mux2_1
X_19138_ _05844_ _05878_ _05879_ _05849_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a22o_1
X_35184_ clknet_leaf_393_CLK _03298_ VGND VGND VPWR VPWR registers\[18\]\[34\] sky130_fd_sc_hd__dfxtp_1
X_32396_ clknet_leaf_166_CLK _00510_ VGND VGND VPWR VPWR registers\[61\]\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34135_ clknet_leaf_106_CLK _02249_ VGND VGND VPWR VPWR registers\[34\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_238_1429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_31347_ _14172_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__clkbuf_1
X_19069_ _05540_ _05810_ _05811_ _05545_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__a22o_1
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21100_ _07783_ _07784_ _07785_ _07786_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__a22o_1
XFILLER_12_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34066_ clknet_leaf_122_CLK _02180_ VGND VGND VPWR VPWR registers\[35\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_22080_ _08469_ _08737_ _08738_ _08472_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__a22o_1
X_31278_ _14136_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33017_ clknet_leaf_285_CLK _01131_ VGND VGND VPWR VPWR registers\[52\]\[43\] sky130_fd_sc_hd__dfxtp_1
X_21031_ _07340_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__clkbuf_4
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30229_ registers\[15\]\[16\] _12968_ _13577_ VGND VGND VPWR VPWR _13584_ sky130_fd_sc_hd__mux2_1
XFILLER_47_1457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_330_CLK clknet_6_45__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_330_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_248_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_234_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25770_ _10760_ registers\[47\]\[14\] _11170_ VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__mux2_1
X_34968_ clknet_leaf_1_CLK _03082_ VGND VGND VPWR VPWR registers\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_22982_ net27 VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24721_ _09510_ registers\[54\]\[0\] _10587_ VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__mux2_1
X_21933_ _08462_ _08594_ _08595_ _08467_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__a22o_1
X_33919_ clknet_leaf_269_CLK _02033_ VGND VGND VPWR VPWR registers\[38\]\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_55_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_853 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34899_ clknet_leaf_101_CLK _03013_ VGND VGND VPWR VPWR registers\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27440_ _11742_ registers\[35\]\[6\] _12078_ VGND VGND VPWR VPWR _12085_ sky130_fd_sc_hd__mux2_1
X_24652_ _10550_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21864_ _08529_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__buf_6
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_215_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23603_ _09963_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
X_20815_ registers\[48\]\[4\] registers\[49\]\[4\] registers\[50\]\[4\] registers\[51\]\[4\]
+ _07319_ _07320_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__mux4_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_1444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24583_ _10513_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_397_CLK clknet_6_32__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_397_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_27371_ _12048_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21795_ _07312_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__buf_2
XFILLER_168_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29110_ net11 VGND VGND VPWR VPWR _12974_ sky130_fd_sc_hd__clkbuf_4
X_23534_ _09926_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26322_ _11442_ VGND VGND VPWR VPWR _11465_ sky130_fd_sc_hd__clkbuf_4
X_20746_ _07366_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__buf_6
XFILLER_243_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29041_ _12927_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__clkbuf_1
X_26253_ _10838_ registers\[44\]\[51\] _11427_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_149_CLK clknet_6_29__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_149_CLK
+ sky130_fd_sc_hd__clkbuf_16
X_23465_ _09552_ registers\[19\]\[18\] _09881_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__mux2_1
X_20677_ registers\[24\]\[0\] registers\[25\]\[0\] registers\[26\]\[0\] registers\[27\]\[0\]
+ _07374_ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__mux4_1
XFILLER_17_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_811 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25204_ _10872_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22416_ _09062_ _09065_ _08759_ VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__o21ba_1
XFILLER_178_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26184_ _11392_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
X_23396_ _09852_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
X_25135_ _10827_ registers\[52\]\[46\] _10815_ VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__mux2_1
X_22347_ _08761_ _08997_ _08998_ _08764_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__a22o_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29943_ _13433_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__clkbuf_1
X_25066_ net17 VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__buf_2
X_22278_ registers\[28\]\[45\] registers\[29\]\[45\] registers\[30\]\[45\] registers\[31\]\[45\]
+ _08835_ _08836_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__mux4_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24017_ _09556_ registers\[5\]\[20\] _10183_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__mux2_1
X_21229_ registers\[36\]\[16\] registers\[37\]\[16\] registers\[38\]\[16\] registers\[39\]\[16\]
+ _07606_ _07607_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__mux4_1
XFILLER_215_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29874_ _13352_ VGND VGND VPWR VPWR _13397_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_321_CLK clknet_6_38__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_321_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_239_918 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28825_ _12814_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28756_ _11841_ registers\[26\]\[53\] _12774_ VGND VGND VPWR VPWR _12778_ sky130_fd_sc_hd__mux2_1
X_16770_ _14546_ VGND VGND VPWR VPWR _15264_ sky130_fd_sc_hd__buf_4
XFILLER_247_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25968_ _10823_ registers\[46\]\[44\] _11274_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__mux2_1
XFILLER_93_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27707_ _12226_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__clkbuf_1
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24919_ _09577_ registers\[53\]\[30\] _10691_ VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__mux2_1
XFILLER_58_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28687_ _11771_ registers\[26\]\[20\] _12741_ VGND VGND VPWR VPWR _12742_ sky130_fd_sc_hd__mux2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25899_ _10754_ registers\[46\]\[11\] _11241_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__mux2_1
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_233_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18440_ registers\[32\]\[2\] registers\[33\]\[2\] registers\[34\]\[2\] registers\[35\]\[2\]
+ _05068_ _05070_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__mux4_1
XFILLER_233_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27638_ registers\[34\]\[35\] _10378_ _12184_ VGND VGND VPWR VPWR _12190_ sky130_fd_sc_hd__mux2_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18371_ _05133_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__buf_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27569_ registers\[34\]\[2\] _10309_ _12151_ VGND VGND VPWR VPWR _12154_ sky130_fd_sc_hd__mux2_1
XFILLER_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_388_CLK clknet_6_34__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_388_CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29308_ _13099_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__clkbuf_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ registers\[24\]\[35\] registers\[25\]\[35\] registers\[26\]\[35\] registers\[27\]\[35\]
+ _15768_ _15769_ VGND VGND VPWR VPWR _15801_ sky130_fd_sc_hd__mux4_1
XFILLER_14_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30580_ _09806_ registers\[13\]\[54\] _13764_ VGND VGND VPWR VPWR _13769_ sky130_fd_sc_hd__mux2_1
XFILLER_18_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29239_ _13061_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17253_ registers\[4\]\[33\] registers\[5\]\[33\] registers\[6\]\[33\] registers\[7\]\[33\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15734_ sky130_fd_sc_hd__mux4_1
XFILLER_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16204_ _14691_ _14698_ _14707_ _14714_ VGND VGND VPWR VPWR _14715_ sky130_fd_sc_hd__or4_2
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32250_ clknet_leaf_281_CLK _00364_ VGND VGND VPWR VPWR registers\[39\]\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17184_ _15487_ _15665_ _15666_ _15490_ VGND VGND VPWR VPWR _15667_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31201_ _14095_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16135_ _14647_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32181_ clknet_leaf_485_CLK _00295_ VGND VGND VPWR VPWR registers\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31132_ registers\[0\]\[60\] _13060_ _13992_ VGND VGND VPWR VPWR _14059_ sky130_fd_sc_hd__mux2_1
X_16066_ registers\[4\]\[0\] registers\[5\]\[0\] registers\[6\]\[0\] registers\[7\]\[0\]
+ _14577_ _14579_ VGND VGND VPWR VPWR _14580_ sky130_fd_sc_hd__mux4_1
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_237_1473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_1023 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_912 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31063_ registers\[0\]\[27\] _12991_ _14015_ VGND VGND VPWR VPWR _14023_ sky130_fd_sc_hd__mux2_1
X_35940_ clknet_leaf_469_CLK _04054_ VGND VGND VPWR VPWR registers\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_312_CLK clknet_6_37__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_312_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30014_ registers\[17\]\[42\] _13023_ _13468_ VGND VGND VPWR VPWR _13471_ sky130_fd_sc_hd__mux2_1
X_19825_ registers\[56\]\[41\] registers\[57\]\[41\] registers\[58\]\[41\] registers\[59\]\[41\]
+ _06301_ _06434_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__mux4_1
X_35871_ clknet_leaf_480_CLK _03985_ VGND VGND VPWR VPWR registers\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_57_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_34822_ clknet_leaf_219_CLK _02936_ VGND VGND VPWR VPWR registers\[24\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19756_ _06476_ _06479_ _06169_ _06170_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__o211a_1
X_16968_ _15453_ _15456_ _15288_ VGND VGND VPWR VPWR _15457_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18707_ _05137_ _05459_ _05460_ _05147_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__a22o_1
XFILLER_133_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34753_ clknet_leaf_224_CLK _02867_ VGND VGND VPWR VPWR registers\[25\]\[51\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_5_16_0_CLK clknet_2_2_0_CLK VGND VGND VPWR VPWR clknet_5_16_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31965_ clknet_leaf_4_CLK _00134_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
X_19687_ _06374_ _06411_ _06412_ _06377_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__a22o_1
X_16899_ registers\[12\]\[23\] registers\[13\]\[23\] registers\[14\]\[23\] registers\[15\]\[23\]
+ _15388_ _15389_ VGND VGND VPWR VPWR _15390_ sky130_fd_sc_hd__mux4_1
X_33704_ clknet_leaf_429_CLK _01818_ VGND VGND VPWR VPWR registers\[41\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_18638_ _05150_ _05392_ _05393_ _05160_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__a22o_1
X_30916_ registers\[10\]\[21\] _12979_ _13944_ VGND VGND VPWR VPWR _13946_ sky130_fd_sc_hd__mux2_1
X_34684_ clknet_leaf_188_CLK _02798_ VGND VGND VPWR VPWR registers\[26\]\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_897 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31896_ _09771_ registers\[49\]\[38\] _14452_ VGND VGND VPWR VPWR _14461_ sky130_fd_sc_hd__mux2_1
XFILLER_224_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33635_ clknet_leaf_55_CLK _01749_ VGND VGND VPWR VPWR registers\[42\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_30847_ _13909_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_240_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18569_ _05323_ _05326_ _05163_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_379_CLK clknet_6_40__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_379_CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_212_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20600_ registers\[44\]\[0\] registers\[45\]\[0\] registers\[46\]\[0\] registers\[47\]\[0\]
+ _07297_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__mux4_1
XFILLER_75_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21580_ _08119_ _08251_ _08252_ _08124_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__a22o_1
X_33566_ clknet_leaf_27_CLK _01680_ VGND VGND VPWR VPWR registers\[43\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_244_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30778_ _13850_ VGND VGND VPWR VPWR _13873_ sky130_fd_sc_hd__buf_4
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_221_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1038 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35305_ clknet_leaf_403_CLK _03419_ VGND VGND VPWR VPWR registers\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_20531_ _05040_ _07230_ _07231_ _05050_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__a22o_1
X_32517_ clknet_leaf_200_CLK _00631_ VGND VGND VPWR VPWR registers\[60\]\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_1188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_33497_ clknet_leaf_31_CLK _01611_ VGND VGND VPWR VPWR registers\[44\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23250_ net28 VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__clkbuf_4
X_35236_ clknet_leaf_447_CLK _03350_ VGND VGND VPWR VPWR registers\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_32448_ clknet_leaf_199_CLK _00562_ VGND VGND VPWR VPWR registers\[29\]\[50\] sky130_fd_sc_hd__dfxtp_1
X_20462_ registers\[56\]\[60\] registers\[57\]\[60\] registers\[58\]\[60\] registers\[59\]\[60\]
+ _06987_ _05152_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__mux4_1
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22201_ registers\[0\]\[43\] registers\[1\]\[43\] registers\[2\]\[43\] registers\[3\]\[43\]
+ _08752_ _08753_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__mux4_1
XFILLER_118_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_203_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23181_ _09720_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_119_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35167_ clknet_leaf_2_CLK _03281_ VGND VGND VPWR VPWR registers\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_20393_ _07077_ _07084_ _07091_ _07098_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__or4_2
X_32379_ clknet_leaf_287_CLK _00493_ VGND VGND VPWR VPWR registers\[61\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34118_ clknet_leaf_248_CLK _02232_ VGND VGND VPWR VPWR registers\[35\]\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22132_ registers\[8\]\[41\] registers\[9\]\[41\] registers\[10\]\[41\] registers\[11\]\[41\]
+ _08577_ _08578_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__mux4_1
XFILLER_238_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput230 net230 VGND VGND VPWR VPWR D3[20] sky130_fd_sc_hd__buf_2
X_35098_ clknet_leaf_10_CLK _03212_ VGND VGND VPWR VPWR registers\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput241 net241 VGND VGND VPWR VPWR D3[30] sky130_fd_sc_hd__buf_2
Xoutput252 net252 VGND VGND VPWR VPWR D3[40] sky130_fd_sc_hd__buf_2
XTAP_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_34049_ clknet_leaf_260_CLK _02163_ VGND VGND VPWR VPWR registers\[36\]\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput263 net263 VGND VGND VPWR VPWR D3[50] sky130_fd_sc_hd__buf_2
X_26940_ net32 VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__clkbuf_4
X_22063_ _08719_ _08722_ _08416_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__o21ba_1
XTAP_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_303_CLK clknet_6_50__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_303_CLK
+ sky130_fd_sc_hd__clkbuf_16
Xoutput274 net274 VGND VGND VPWR VPWR D3[60] sky130_fd_sc_hd__buf_2
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_248_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_21014_ registers\[40\]\[10\] registers\[41\]\[10\] registers\[42\]\[10\] registers\[43\]\[10\]
+ _07434_ _07435_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__mux4_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26871_ _11762_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__clkbuf_1
XTAP_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_28610_ _11830_ registers\[27\]\[48\] _12692_ VGND VGND VPWR VPWR _12701_ sky130_fd_sc_hd__mux2_1
X_25822_ _10812_ registers\[47\]\[39\] _11192_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__mux2_1
XFILLER_229_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29590_ registers\[20\]\[33\] _13004_ _13244_ VGND VGND VPWR VPWR _13248_ sky130_fd_sc_hd__mux2_1
XFILLER_216_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_28541_ _11761_ registers\[27\]\[15\] _12659_ VGND VGND VPWR VPWR _12665_ sky130_fd_sc_hd__mux2_1
X_25753_ _10743_ registers\[47\]\[6\] _11159_ VGND VGND VPWR VPWR _11166_ sky130_fd_sc_hd__mux2_1
XFILLER_244_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22965_ _09572_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_243_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_228_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_24704_ _10577_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_812 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28472_ _12628_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__clkbuf_1
X_21916_ registers\[0\]\[35\] registers\[1\]\[35\] registers\[2\]\[35\] registers\[3\]\[35\]
+ _08409_ _08410_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__mux4_1
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22896_ _09525_ registers\[62\]\[5\] _09515_ VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__mux2_1
X_25684_ _11128_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27423_ _12075_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_215_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21847_ registers\[8\]\[33\] registers\[9\]\[33\] registers\[10\]\[33\] registers\[11\]\[33\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__mux4_1
X_24635_ _10541_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__clkbuf_1
X_24566_ _10503_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27354_ _12039_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__clkbuf_1
X_21778_ _08442_ _08445_ _08405_ _08406_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__o211a_1
XFILLER_168_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26305_ _11456_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
X_20729_ _07373_ _07425_ _07426_ _07383_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__a22o_1
XFILLER_156_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23517_ _09917_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
X_27285_ _11857_ registers\[37\]\[61\] _11935_ VGND VGND VPWR VPWR _12003_ sky130_fd_sc_hd__mux2_1
X_24497_ _10467_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_29024_ registers\[24\]\[52\] _10414_ _12916_ VGND VGND VPWR VPWR _12919_ sky130_fd_sc_hd__mux2_1
XFILLER_17_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_26236_ _10821_ registers\[44\]\[43\] _11416_ VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__mux2_1
X_23448_ _09869_ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__buf_4
XFILLER_104_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23379_ _09843_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
X_26167_ _10751_ registers\[44\]\[10\] _11383_ VGND VGND VPWR VPWR _11384_ sky130_fd_sc_hd__mux2_1
X_25118_ _10816_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26098_ _11347_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17940_ registers\[32\]\[53\] registers\[33\]\[53\] registers\[34\]\[53\] registers\[35\]\[53\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__mux4_1
X_29926_ registers\[17\]\[0\] _12931_ _13424_ VGND VGND VPWR VPWR _13425_ sky130_fd_sc_hd__mux2_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_25049_ _10769_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17871_ registers\[40\]\[51\] registers\[41\]\[51\] registers\[42\]\[51\] registers\[43\]\[51\]
+ _04334_ _04335_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__mux4_1
XFILLER_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29857_ _13388_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19610_ registers\[52\]\[35\] registers\[53\]\[35\] registers\[54\]\[35\] registers\[55\]\[35\]
+ _06026_ _06027_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__mux4_1
XFILLER_120_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16822_ registers\[60\]\[21\] registers\[61\]\[21\] registers\[62\]\[21\] registers\[63\]\[21\]
+ _15070_ _15207_ VGND VGND VPWR VPWR _15315_ sky130_fd_sc_hd__mux4_1
X_28808_ _12805_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29788_ _13351_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19541_ registers\[48\]\[33\] registers\[49\]\[33\] registers\[50\]\[33\] registers\[51\]\[33\]
+ _06093_ _06094_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux4_1
XFILLER_235_921 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_219_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_28739_ _11824_ registers\[26\]\[45\] _12763_ VGND VGND VPWR VPWR _12769_ sky130_fd_sc_hd__mux2_1
X_16753_ _15139_ _15246_ _15247_ _15142_ VGND VGND VPWR VPWR _15248_ sky130_fd_sc_hd__a22o_1
XFILLER_98_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31750_ _14384_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__clkbuf_1
X_19472_ registers\[56\]\[31\] registers\[57\]\[31\] registers\[58\]\[31\] registers\[59\]\[31\]
+ _05958_ _06091_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__mux4_1
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16684_ _15144_ _15179_ _15180_ _15147_ VGND VGND VPWR VPWR _15181_ sky130_fd_sc_hd__a22o_1
XFILLER_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18423_ registers\[12\]\[1\] registers\[13\]\[1\] registers\[14\]\[1\] registers\[15\]\[1\]
+ _05121_ _05123_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__mux4_1
XFILLER_179_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30701_ _13832_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31681_ _14347_ VGND VGND VPWR VPWR _14348_ sky130_fd_sc_hd__buf_4
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_33420_ clknet_leaf_164_CLK _01534_ VGND VGND VPWR VPWR registers\[46\]\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__buf_4
XFILLER_159_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30632_ _13796_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _15780_ _15783_ _15612_ VGND VGND VPWR VPWR _15784_ sky130_fd_sc_hd__o21ba_1
X_33351_ clknet_leaf_250_CLK _01465_ VGND VGND VPWR VPWR registers\[47\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18285_ net79 net80 VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nor2_4
XFILLER_159_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30563_ _09788_ registers\[13\]\[46\] _13753_ VGND VGND VPWR VPWR _13760_ sky130_fd_sc_hd__mux2_1
X_32302_ clknet_leaf_394_CLK _00416_ VGND VGND VPWR VPWR registers\[19\]\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17236_ registers\[44\]\[33\] registers\[45\]\[33\] registers\[46\]\[33\] registers\[47\]\[33\]
+ _15607_ _15608_ VGND VGND VPWR VPWR _15717_ sky130_fd_sc_hd__mux4_1
X_36070_ clknet_leaf_439_CLK _04184_ VGND VGND VPWR VPWR registers\[59\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_33282_ clknet_leaf_259_CLK _01396_ VGND VGND VPWR VPWR registers\[48\]\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1071 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_30494_ _09685_ registers\[13\]\[13\] _13720_ VGND VGND VPWR VPWR _13724_ sky130_fd_sc_hd__mux2_1
XFILLER_174_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35021_ clknet_leaf_145_CLK _03135_ VGND VGND VPWR VPWR registers\[21\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_32233_ clknet_leaf_146_CLK _00347_ VGND VGND VPWR VPWR registers\[9\]\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_17167_ _15334_ _15648_ _15649_ _15339_ VGND VGND VPWR VPWR _15650_ sky130_fd_sc_hd__a22o_1
XFILLER_116_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16118_ _14540_ _14629_ _14630_ _14551_ VGND VGND VPWR VPWR _14631_ sky130_fd_sc_hd__a22o_1
X_32164_ clknet_leaf_108_CLK _00278_ VGND VGND VPWR VPWR registers\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17098_ registers\[48\]\[29\] registers\[49\]\[29\] registers\[50\]\[29\] registers\[51\]\[29\]
+ _15544_ _15545_ VGND VGND VPWR VPWR _15583_ sky130_fd_sc_hd__mux4_1
XFILLER_171_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31115_ _14050_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16049_ _14562_ VGND VGND VPWR VPWR _14563_ sky130_fd_sc_hd__buf_6
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_32095_ clknet_leaf_485_CLK _00008_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dfxtp_1
XFILLER_130_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35923_ clknet_leaf_77_CLK _04037_ VGND VGND VPWR VPWR registers\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31046_ registers\[0\]\[19\] _12974_ _14004_ VGND VGND VPWR VPWR _14014_ sky130_fd_sc_hd__mux2_1
XFILLER_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19808_ registers\[28\]\[40\] registers\[29\]\[40\] registers\[30\]\[40\] registers\[31\]\[40\]
+ _06256_ _06257_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__mux4_1
X_35854_ clknet_leaf_108_CLK _03968_ VGND VGND VPWR VPWR registers\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_245_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_34805_ clknet_leaf_414_CLK _02919_ VGND VGND VPWR VPWR registers\[24\]\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19739_ _06432_ _06447_ _06456_ _06463_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__or4_2
X_35785_ clknet_leaf_216_CLK _03899_ VGND VGND VPWR VPWR registers\[0\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_32997_ clknet_leaf_438_CLK _01111_ VGND VGND VPWR VPWR registers\[52\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_231_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22750_ registers\[20\]\[59\] registers\[21\]\[59\] registers\[22\]\[59\] registers\[23\]\[59\]
+ _09111_ _09112_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__mux4_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31948_ _09825_ registers\[49\]\[63\] _14418_ VGND VGND VPWR VPWR _14488_ sky130_fd_sc_hd__mux2_1
X_34736_ clknet_leaf_411_CLK _02850_ VGND VGND VPWR VPWR registers\[25\]\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_21701_ registers\[52\]\[29\] registers\[53\]\[29\] registers\[54\]\[29\] registers\[55\]\[29\]
+ _08262_ _08263_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__mux4_1
X_22681_ _07276_ _09321_ _09322_ _07286_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__a22o_1
X_34667_ clknet_leaf_452_CLK _02781_ VGND VGND VPWR VPWR registers\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31879_ _14418_ VGND VGND VPWR VPWR _14452_ sky130_fd_sc_hd__buf_4
X_24420_ registers\[57\]\[56\] _10422_ _10410_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__mux2_1
X_33618_ clknet_leaf_125_CLK _01732_ VGND VGND VPWR VPWR registers\[42\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_21632_ registers\[8\]\[27\] registers\[9\]\[27\] registers\[10\]\[27\] registers\[11\]\[27\]
+ _08234_ _08235_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__mux4_1
XFILLER_178_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34598_ clknet_leaf_450_CLK _02712_ VGND VGND VPWR VPWR registers\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_240_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24351_ net28 VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__buf_4
XFILLER_51_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33549_ clknet_leaf_172_CLK _01663_ VGND VGND VPWR VPWR registers\[44\]\[63\] sky130_fd_sc_hd__dfxtp_1
X_21563_ registers\[0\]\[25\] registers\[1\]\[25\] registers\[2\]\[25\] registers\[3\]\[25\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__mux4_1
XFILLER_205_1269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23302_ _09796_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__clkbuf_1
X_20514_ _07215_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__buf_4
X_27070_ _11890_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_1
X_24282_ _10329_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_909 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_21494_ registers\[8\]\[23\] registers\[9\]\[23\] registers\[10\]\[23\] registers\[11\]\[23\]
+ _07891_ _07892_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__mux4_1
X_26021_ _10741_ registers\[45\]\[5\] _11301_ VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__mux2_1
X_35219_ clknet_leaf_102_CLK _03333_ VGND VGND VPWR VPWR registers\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_23233_ _09750_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
X_20445_ _07145_ _07148_ _06866_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__o21ba_1
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36199_ clknet_leaf_98_CLK _00081_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_CLK clknet_6_19__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_80_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23164_ _09711_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
X_20376_ registers\[52\]\[57\] registers\[53\]\[57\] registers\[54\]\[57\] registers\[55\]\[57\]
+ _05043_ _05046_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__mux4_1
XTAP_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22115_ _08765_ _08772_ _08773_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__o21ba_1
XTAP_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23095_ _09663_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_216_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27972_ _11732_ registers\[31\]\[1\] _12364_ VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__mux2_1
XFILLER_175_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_248_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_29711_ _13311_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26923_ _11797_ registers\[3\]\[32\] _11793_ VGND VGND VPWR VPWR _11798_ sky130_fd_sc_hd__mux2_1
X_22046_ registers\[44\]\[39\] registers\[45\]\[39\] registers\[46\]\[39\] registers\[47\]\[39\]
+ _08392_ _08393_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__mux4_1
XTAP_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_1387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_248_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_212_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29642_ registers\[20\]\[58\] _13056_ _13266_ VGND VGND VPWR VPWR _13275_ sky130_fd_sc_hd__mux2_1
XTAP_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26854_ _11729_ VGND VGND VPWR VPWR _11751_ sky130_fd_sc_hd__buf_4
XFILLER_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_937 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_1382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25805_ _11193_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29573_ registers\[20\]\[25\] _12987_ _13233_ VGND VGND VPWR VPWR _13239_ sky130_fd_sc_hd__mux2_1
X_26785_ _11709_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_23997_ _10173_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
X_28524_ _11744_ registers\[27\]\[7\] _12648_ VGND VGND VPWR VPWR _12656_ sky130_fd_sc_hd__mux2_1
XFILLER_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25736_ _11155_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_22948_ net15 VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__buf_2
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28455_ _12619_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_216_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25667_ registers\[48\]\[30\] _10367_ _11119_ VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__mux2_1
X_22879_ _09513_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__buf_12
XFILLER_44_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27406_ registers\[36\]\[54\] _10418_ _12062_ VGND VGND VPWR VPWR _12067_ sky130_fd_sc_hd__mux2_1
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_227_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24618_ _10532_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
X_28386_ _12583_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__clkbuf_1
X_25598_ _11081_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_883 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_27337_ registers\[36\]\[21\] _10349_ _12029_ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__mux2_1
XFILLER_184_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24549_ _10494_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_169_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18070_ _04683_ _04838_ _04839_ _04686_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a22o_1
X_27268_ _11994_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_29007_ registers\[24\]\[44\] _10397_ _12905_ VGND VGND VPWR VPWR _12910_ sky130_fd_sc_hd__mux2_1
X_17021_ _14573_ VGND VGND VPWR VPWR _15508_ sky130_fd_sc_hd__clkbuf_8
XFILLER_172_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26219_ _10804_ registers\[44\]\[35\] _11405_ VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__mux2_1
X_27199_ _11935_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_71_CLK clknet_6_24__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_71_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18972_ registers\[56\]\[17\] registers\[57\]\[17\] registers\[58\]\[17\] registers\[59\]\[17\]
+ _05615_ _05405_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__mux4_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1700 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1711 _00164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17923_ _04481_ _04696_ _04697_ _04484_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a22o_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29909_ _13415_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1722 _00169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1733 _00178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1744 _05049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1755 _07303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32920_ clknet_leaf_66_CLK _01034_ VGND VGND VPWR VPWR registers\[53\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1766 _08407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17854_ _04626_ _04629_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__o21ba_1
XFILLER_121_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1777 _11935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1788 _14571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_227_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16805_ registers\[20\]\[20\] registers\[21\]\[20\] registers\[22\]\[20\] registers\[23\]\[20\]
+ _15297_ _15298_ VGND VGND VPWR VPWR _15299_ sky130_fd_sc_hd__mux4_1
X_32851_ clknet_leaf_181_CLK _00965_ VGND VGND VPWR VPWR registers\[54\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_17785_ registers\[24\]\[48\] registers\[25\]\[48\] registers\[26\]\[48\] registers\[27\]\[48\]
+ _04424_ _04425_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__mux4_1
XFILLER_43_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31802_ _14411_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__clkbuf_1
X_19524_ _06182_ _06253_ _06254_ _06185_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__a22o_1
X_35570_ clknet_leaf_380_CLK _03684_ VGND VGND VPWR VPWR registers\[12\]\[36\] sky130_fd_sc_hd__dfxtp_1
X_16736_ _14518_ VGND VGND VPWR VPWR _15231_ sky130_fd_sc_hd__buf_4
XFILLER_228_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32782_ clknet_leaf_179_CLK _00896_ VGND VGND VPWR VPWR registers\[55\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_34521_ clknet_leaf_21_CLK _02635_ VGND VGND VPWR VPWR registers\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_19455_ registers\[28\]\[30\] registers\[29\]\[30\] registers\[30\]\[30\] registers\[31\]\[30\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__mux4_1
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31733_ _14375_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16667_ _14571_ VGND VGND VPWR VPWR _15164_ sky130_fd_sc_hd__buf_4
X_18406_ _05040_ _05166_ _05167_ _05050_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a22o_1
XFILLER_90_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34452_ clknet_leaf_88_CLK _02566_ VGND VGND VPWR VPWR registers\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_31664_ registers\[63\]\[56\] net52 _14332_ VGND VGND VPWR VPWR _14339_ sky130_fd_sc_hd__mux2_1
XFILLER_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19386_ _06089_ _06104_ _06113_ _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__or4_4
X_16598_ _14998_ _15095_ _15096_ _15001_ VGND VGND VPWR VPWR _15097_ sky130_fd_sc_hd__a22o_1
X_33403_ clknet_leaf_278_CLK _01517_ VGND VGND VPWR VPWR registers\[46\]\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30615_ _13787_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__clkbuf_1
X_18337_ _05065_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__clkbuf_4
X_34383_ clknet_leaf_111_CLK _02497_ VGND VGND VPWR VPWR registers\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_31595_ registers\[63\]\[23\] net16 _14299_ VGND VGND VPWR VPWR _14303_ sky130_fd_sc_hd__mux2_1
XFILLER_241_1469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_36122_ clknet_leaf_52_CLK _04236_ VGND VGND VPWR VPWR registers\[49\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33334_ clknet_leaf_341_CLK _01448_ VGND VGND VPWR VPWR registers\[47\]\[40\] sky130_fd_sc_hd__dfxtp_1
X_18268_ _14558_ _05030_ _05031_ _14568_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__a22o_1
X_30546_ _09771_ registers\[13\]\[38\] _13742_ VGND VGND VPWR VPWR _13751_ sky130_fd_sc_hd__mux2_1
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36053_ clknet_leaf_64_CLK _04167_ VGND VGND VPWR VPWR registers\[59\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_17219_ registers\[4\]\[32\] registers\[5\]\[32\] registers\[6\]\[32\] registers\[7\]\[32\]
+ _15560_ _15561_ VGND VGND VPWR VPWR _15701_ sky130_fd_sc_hd__mux4_1
XFILLER_162_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33265_ clknet_leaf_366_CLK _01379_ VGND VGND VPWR VPWR registers\[48\]\[35\] sky130_fd_sc_hd__dfxtp_1
X_18199_ registers\[8\]\[61\] registers\[9\]\[61\] registers\[10\]\[61\] registers\[11\]\[61\]
+ _14503_ _14505_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__mux4_1
X_30477_ _09668_ registers\[13\]\[5\] _13709_ VGND VGND VPWR VPWR _13715_ sky130_fd_sc_hd__mux2_1
XFILLER_144_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_CLK clknet_6_26__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_62_CLK sky130_fd_sc_hd__clkbuf_16
X_35004_ clknet_leaf_307_CLK _03118_ VGND VGND VPWR VPWR registers\[21\]\[46\] sky130_fd_sc_hd__dfxtp_1
X_20230_ _06868_ _06939_ _06940_ _06871_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__a22o_1
X_32216_ clknet_leaf_288_CLK _00330_ VGND VGND VPWR VPWR registers\[9\]\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33196_ clknet_leaf_390_CLK _01310_ VGND VGND VPWR VPWR registers\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32147_ clknet_leaf_119_CLK _00261_ VGND VGND VPWR VPWR registers\[39\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_20161_ registers\[28\]\[50\] registers\[29\]\[50\] registers\[30\]\[50\] registers\[31\]\[50\]
+ _06599_ _06600_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__mux4_1
XFILLER_157_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20092_ _06775_ _06790_ _06799_ _06806_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__or4_4
X_32078_ clknet_leaf_491_CLK _00000_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35906_ clknet_leaf_264_CLK _04020_ VGND VGND VPWR VPWR registers\[7\]\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_31029_ _14005_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__clkbuf_1
X_23920_ _09596_ registers\[60\]\[39\] _10122_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__mux2_1
XFILLER_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_35837_ clknet_leaf_288_CLK _03951_ VGND VGND VPWR VPWR registers\[8\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_23851_ _09527_ registers\[60\]\[6\] _10089_ VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__mux2_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_242_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_22802_ registers\[12\]\[61\] registers\[13\]\[61\] registers\[14\]\[61\] registers\[15\]\[61\]
+ _09202_ _09203_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__mux4_1
XFILLER_66_981 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26570_ _10749_ registers\[41\]\[9\] _11586_ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__mux2_1
XANTENNA_608 _05111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ registers\[60\]\[9\] registers\[61\]\[9\] registers\[62\]\[9\] registers\[63\]\[9\]
+ _07512_ _07649_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__mux4_1
XANTENNA_619 _05116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35768_ clknet_leaf_316_CLK _03882_ VGND VGND VPWR VPWR registers\[0\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_23782_ _09594_ registers\[29\]\[38\] _10050_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__mux2_1
XFILLER_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25521_ _11041_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22733_ registers\[48\]\[59\] registers\[49\]\[59\] registers\[50\]\[59\] registers\[51\]\[59\]
+ _07327_ _07392_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__mux4_1
XFILLER_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34719_ clknet_leaf_9_CLK _02833_ VGND VGND VPWR VPWR registers\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_246_1358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_35699_ clknet_leaf_383_CLK _03813_ VGND VGND VPWR VPWR registers\[10\]\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28240_ registers\[2\]\[0\] _10303_ _12506_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__mux2_1
X_22664_ _09306_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
X_25452_ _10856_ registers\[50\]\[60\] _10936_ VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__mux2_1
XFILLER_240_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_205_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24403_ _10411_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
X_21615_ _08287_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28171_ _12470_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_244_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22595_ _07349_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__buf_4
XFILLER_187_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25383_ _10787_ registers\[50\]\[27\] _10959_ VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__mux2_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27122_ _11917_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__clkbuf_1
X_24334_ _10364_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
X_21546_ registers\[40\]\[25\] registers\[41\]\[25\] registers\[42\]\[25\] registers\[43\]\[25\]
+ _08120_ _08121_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__mux4_1
XFILLER_166_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24265_ registers\[57\]\[6\] _10317_ _10305_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__mux2_1
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27053_ _11881_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_1
X_21477_ _08148_ _08153_ _08087_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__o21ba_1
XFILLER_140_1080 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_CLK clknet_6_13__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_53_CLK sky130_fd_sc_hd__clkbuf_16
X_26004_ _11297_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
X_23216_ _09739_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
X_20428_ registers\[44\]\[59\] registers\[45\]\[59\] registers\[46\]\[59\] registers\[47\]\[59\]
+ _06842_ _06843_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__mux4_1
XFILLER_153_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_953 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24196_ _10278_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23147_ _09698_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20359_ registers\[28\]\[56\] registers\[29\]\[56\] registers\[30\]\[56\] registers\[31\]\[56\]
+ _06942_ _06943_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__mux4_1
XTAP_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1007 _11845_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_1149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1018 _12363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27955_ _12356_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__clkbuf_1
X_23078_ net87 VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__buf_4
XTAP_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1029 _12934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_216_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26906_ net20 VGND VGND VPWR VPWR _11786_ sky130_fd_sc_hd__clkbuf_4
X_22029_ registers\[4\]\[38\] registers\[5\]\[38\] registers\[6\]\[38\] registers\[7\]\[38\]
+ _08688_ _08689_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__mux4_1
XTAP_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27886_ _12320_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29625_ _13210_ VGND VGND VPWR VPWR _13266_ sky130_fd_sc_hd__buf_4
XTAP_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26837_ _11739_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _15825_ _04353_ _04354_ _15828_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a22o_1
X_29556_ registers\[20\]\[17\] _12970_ _13222_ VGND VGND VPWR VPWR _13230_ sky130_fd_sc_hd__mux2_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26768_ _11700_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28507_ _12646_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__clkbuf_1
X_16521_ registers\[28\]\[12\] registers\[29\]\[12\] registers\[30\]\[12\] registers\[31\]\[12\]
+ _15021_ _15022_ VGND VGND VPWR VPWR _15023_ sky130_fd_sc_hd__mux4_1
XFILLER_95_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25719_ registers\[48\]\[55\] _10420_ _11141_ VGND VGND VPWR VPWR _11147_ sky130_fd_sc_hd__mux2_1
XFILLER_216_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_29487_ _13193_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26699_ _11664_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_225_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19240_ registers\[28\]\[24\] registers\[29\]\[24\] registers\[30\]\[24\] registers\[31\]\[24\]
+ _05913_ _05914_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__mux4_1
X_16452_ registers\[20\]\[10\] registers\[21\]\[10\] registers\[22\]\[10\] registers\[23\]\[10\]
+ _14954_ _14955_ VGND VGND VPWR VPWR _14956_ sky130_fd_sc_hd__mux4_1
X_28438_ _11792_ registers\[28\]\[30\] _12610_ VGND VGND VPWR VPWR _12611_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_1442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_231_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19171_ _05839_ _05910_ _05911_ _05842_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__a22o_1
X_28369_ registers\[2\]\[62\] _10434_ _12505_ VGND VGND VPWR VPWR _12574_ sky130_fd_sc_hd__mux2_1
XFILLER_231_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16383_ _14518_ VGND VGND VPWR VPWR _14888_ sky130_fd_sc_hd__buf_6
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18122_ _04887_ _04890_ _04644_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o21ba_1
X_30400_ _13674_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__clkbuf_1
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_223_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31380_ _14189_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_223_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_864 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18053_ registers\[4\]\[56\] registers\[5\]\[56\] registers\[6\]\[56\] registers\[7\]\[56\]
+ _04559_ _04560_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__mux4_1
X_30331_ _13637_ VGND VGND VPWR VPWR _13638_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_44_CLK clknet_6_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_44_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17004_ _15486_ _15491_ _15288_ VGND VGND VPWR VPWR _15492_ sky130_fd_sc_hd__o21ba_1
XANTENNA_4 _00025_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33050_ clknet_leaf_52_CLK _01164_ VGND VGND VPWR VPWR registers\[51\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_30262_ _13601_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__clkbuf_1
X_32001_ clknet_leaf_27_CLK _00174_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_30193_ _13564_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18955_ registers\[16\]\[16\] registers\[17\]\[16\] registers\[18\]\[16\] registers\[19\]\[16\]
+ _05700_ _05701_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__mux4_1
XANTENNA_1530 _09215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_234_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1541 _09793_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1552 _11371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_230_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17906_ _14500_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__clkbuf_8
XFILLER_140_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18886_ _05496_ _05633_ _05634_ _05499_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a22o_1
XANTENNA_1563 _11761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33952_ clknet_leaf_16_CLK _02066_ VGND VGND VPWR VPWR registers\[37\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1574 _13210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1585 _14490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1596 _14548_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ registers\[48\]\[50\] registers\[49\]\[50\] registers\[50\]\[50\] registers\[51\]\[50\]
+ _04543_ _04544_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__mux4_1
X_32903_ clknet_leaf_194_CLK _01017_ VGND VGND VPWR VPWR registers\[54\]\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33883_ clknet_leaf_24_CLK _01997_ VGND VGND VPWR VPWR registers\[38\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_227_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32834_ clknet_leaf_266_CLK _00948_ VGND VGND VPWR VPWR registers\[55\]\[52\] sky130_fd_sc_hd__dfxtp_1
X_35622_ clknet_leaf_465_CLK _03736_ VGND VGND VPWR VPWR registers\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_17768_ _04540_ _04542_ _04545_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a22o_1
XFILLER_212_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1009 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_242_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16719_ _15139_ _15213_ _15214_ _15142_ VGND VGND VPWR VPWR _15215_ sky130_fd_sc_hd__a22o_1
X_19507_ _06232_ _06237_ _06161_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__o21ba_1
X_32765_ clknet_leaf_289_CLK _00879_ VGND VGND VPWR VPWR registers\[56\]\[47\] sky130_fd_sc_hd__dfxtp_1
X_35553_ clknet_leaf_482_CLK _03667_ VGND VGND VPWR VPWR registers\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17699_ _04474_ _04479_ _15963_ _15964_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__o211a_1
Xclkbuf_6_56__f_CLK clknet_5_28_0_CLK VGND VGND VPWR VPWR clknet_6_56__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34504_ clknet_leaf_154_CLK _02618_ VGND VGND VPWR VPWR registers\[2\]\[58\] sky130_fd_sc_hd__dfxtp_1
X_19438_ _06165_ _06168_ _06169_ _06170_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__o211a_1
X_31716_ _14366_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_35484_ clknet_leaf_477_CLK _03598_ VGND VGND VPWR VPWR registers\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_222_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_32696_ clknet_leaf_334_CLK _00810_ VGND VGND VPWR VPWR registers\[57\]\[42\] sky130_fd_sc_hd__dfxtp_1
X_34435_ clknet_leaf_205_CLK _02549_ VGND VGND VPWR VPWR registers\[30\]\[53\] sky130_fd_sc_hd__dfxtp_1
X_31647_ registers\[63\]\[48\] net43 _14321_ VGND VGND VPWR VPWR _14330_ sky130_fd_sc_hd__mux2_1
X_19369_ _06097_ _06103_ _05826_ _05827_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__o211a_1
XFILLER_241_1233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21400_ _08075_ _08076_ _08077_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__a22o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22380_ _07361_ VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__buf_6
X_34366_ clknet_leaf_182_CLK _02480_ VGND VGND VPWR VPWR registers\[31\]\[48\] sky130_fd_sc_hd__dfxtp_1
X_31578_ registers\[63\]\[15\] net7 _14288_ VGND VGND VPWR VPWR _14294_ sky130_fd_sc_hd__mux2_1
XFILLER_157_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_36105_ clknet_leaf_161_CLK _04219_ VGND VGND VPWR VPWR registers\[59\]\[59\] sky130_fd_sc_hd__dfxtp_1
X_33317_ clknet_leaf_59_CLK _01431_ VGND VGND VPWR VPWR registers\[47\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_21331_ _07737_ _08010_ _08011_ _07742_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__a22o_1
XFILLER_11_1201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30529_ _13708_ VGND VGND VPWR VPWR _13742_ sky130_fd_sc_hd__buf_6
XFILLER_191_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_920 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_34297_ clknet_leaf_340_CLK _02411_ VGND VGND VPWR VPWR registers\[32\]\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_CLK clknet_6_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_35_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24050_ _09590_ registers\[5\]\[36\] _10194_ VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__mux2_1
XFILLER_191_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_36036_ clknet_leaf_201_CLK _04150_ VGND VGND VPWR VPWR registers\[63\]\[54\] sky130_fd_sc_hd__dfxtp_1
X_21262_ _07944_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_33248_ clknet_leaf_42_CLK _01362_ VGND VGND VPWR VPWR registers\[48\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_901 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_23001_ _09596_ registers\[62\]\[39\] _09578_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__mux2_1
X_20213_ _06918_ _06923_ _06847_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__o21ba_1
XFILLER_190_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_1289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_33179_ clknet_leaf_476_CLK _01293_ VGND VGND VPWR VPWR registers\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21193_ registers\[40\]\[15\] registers\[41\]\[15\] registers\[42\]\[15\] registers\[43\]\[15\]
+ _07777_ _07778_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__mux4_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_20144_ _06851_ _06854_ _06855_ _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__o211a_1
XFILLER_89_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_213_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27740_ _12243_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__clkbuf_1
X_20075_ _06783_ _06789_ _06512_ _06513_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__o211a_1
X_24952_ _09611_ registers\[53\]\[46\] _10702_ VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__mux2_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_23903_ _10123_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
X_27671_ _12207_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__clkbuf_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_24883_ _09542_ registers\[53\]\[13\] _10669_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__mux2_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29410_ _13153_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_26622_ _11623_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__clkbuf_1
X_23834_ _09646_ registers\[29\]\[63\] _10016_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__mux2_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _00098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_416 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29341_ _09782_ registers\[22\]\[43\] _13113_ VGND VGND VPWR VPWR _13117_ sky130_fd_sc_hd__mux2_1
XANTENNA_427 _00128_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26553_ _11587_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_438 _00139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ registers\[20\]\[8\] registers\[21\]\[8\] registers\[22\]\[8\] registers\[23\]\[8\]
+ _07391_ _07393_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__mux4_1
X_23765_ _10016_ VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__buf_4
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_449 _00160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25504_ _11032_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__clkbuf_1
X_22716_ registers\[24\]\[58\] registers\[25\]\[58\] registers\[26\]\[58\] registers\[27\]\[58\]
+ _09239_ _09240_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__mux4_1
XFILLER_199_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29272_ _09678_ registers\[22\]\[10\] _13080_ VGND VGND VPWR VPWR _13081_ sky130_fd_sc_hd__mux2_1
XFILLER_53_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26484_ _11550_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__clkbuf_1
X_23696_ registers\[61\]\[63\] _09825_ _09942_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__mux2_1
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_241_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_28223_ _12497_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_25435_ _10994_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22647_ _09020_ _09288_ _09289_ _09024_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__a22o_1
XFILLER_224_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_220_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_881 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_28154_ _12461_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__clkbuf_1
X_22578_ _07314_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__buf_6
X_25366_ _10770_ registers\[50\]\[19\] _10948_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__mux2_1
XFILLER_21_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27105_ _11908_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24317_ net16 VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__clkbuf_4
X_28085_ _11845_ registers\[31\]\[55\] _12419_ VGND VGND VPWR VPWR _12425_ sky130_fd_sc_hd__mux2_1
XFILLER_182_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21529_ registers\[0\]\[24\] registers\[1\]\[24\] registers\[2\]\[24\] registers\[3\]\[24\]
+ _08066_ _08067_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__mux4_1
X_25297_ _10921_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_CLK clknet_6_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_26_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27036_ _11872_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24248_ _10306_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_997 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_24179_ _10269_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_28987_ _12899_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__clkbuf_1
XTAP_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net96 VGND VGND VPWR VPWR D1[15] sky130_fd_sc_hd__buf_2
XFILLER_89_870 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18740_ _05350_ _05491_ _05492_ _05353_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__a22o_1
XTAP_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27938_ _12347_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__clkbuf_1
XTAP_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _05350_ _05422_ _05425_ _05353_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__a22o_1
XTAP_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_27869_ _12311_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_248_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ registers\[36\]\[44\] registers\[37\]\[44\] registers\[38\]\[44\] registers\[39\]\[44\]
+ _15850_ _15851_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__mux4_1
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_29608_ _13257_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__clkbuf_1
X_30880_ registers\[10\]\[4\] _12943_ _13922_ VGND VGND VPWR VPWR _13927_ sky130_fd_sc_hd__mux2_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _14500_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__clkbuf_4
X_29539_ registers\[20\]\[9\] _12953_ _13211_ VGND VGND VPWR VPWR _13221_ sky130_fd_sc_hd__mux2_1
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_229_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_950 _10428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16504_ _14855_ _15004_ _15005_ _14861_ VGND VGND VPWR VPWR _15006_ sky130_fd_sc_hd__a22o_1
XFILLER_60_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_961 _10848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32550_ clknet_leaf_456_CLK _00664_ VGND VGND VPWR VPWR registers\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_204_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_972 _11085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17484_ registers\[48\]\[40\] registers\[49\]\[40\] registers\[50\]\[40\] registers\[51\]\[40\]
+ _15887_ _15888_ VGND VGND VPWR VPWR _15958_ sky130_fd_sc_hd__mux4_1
XFILLER_220_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_983 _11371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_994 _11761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_31501_ _14253_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__clkbuf_1
X_19223_ _05090_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__buf_8
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_16435_ _14564_ VGND VGND VPWR VPWR _14939_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_32481_ clknet_leaf_444_CLK _00595_ VGND VGND VPWR VPWR registers\[60\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34220_ clknet_leaf_322_CLK _02334_ VGND VGND VPWR VPWR registers\[33\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31432_ _14205_ VGND VGND VPWR VPWR _14217_ sky130_fd_sc_hd__buf_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19154_ _05889_ _05894_ _05818_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__o21ba_1
XFILLER_201_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16366_ _14796_ _14870_ _14871_ _14799_ VGND VGND VPWR VPWR _14872_ sky130_fd_sc_hd__a22o_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18105_ registers\[60\]\[58\] registers\[61\]\[58\] registers\[62\]\[58\] registers\[63\]\[58\]
+ _04755_ _14594_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__mux4_1
XFILLER_125_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_34151_ clknet_leaf_431_CLK _02265_ VGND VGND VPWR VPWR registers\[34\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_19085_ _05822_ _05825_ _05826_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o211a_1
X_31363_ registers\[7\]\[41\] net36 _14179_ VGND VGND VPWR VPWR _14181_ sky130_fd_sc_hd__mux2_1
X_16297_ _14801_ _14802_ _14803_ _14804_ VGND VGND VPWR VPWR _14805_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_CLK clknet_6_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_17_CLK sky130_fd_sc_hd__clkbuf_16
X_33102_ clknet_leaf_74_CLK _01216_ VGND VGND VPWR VPWR registers\[50\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_18036_ registers\[32\]\[56\] registers\[33\]\[56\] registers\[34\]\[56\] registers\[35\]\[56\]
+ _04573_ _04574_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__mux4_1
X_30314_ _13628_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_34082_ clknet_leaf_46_CLK _02196_ VGND VGND VPWR VPWR registers\[35\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_31294_ _14144_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33033_ clknet_leaf_193_CLK _01147_ VGND VGND VPWR VPWR registers\[52\]\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_30245_ _13592_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1005 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_30176_ registers\[16\]\[55\] _13050_ _13550_ VGND VGND VPWR VPWR _13556_ sky130_fd_sc_hd__mux2_1
X_19987_ registers\[44\]\[46\] registers\[45\]\[46\] registers\[46\]\[46\] registers\[47\]\[46\]
+ _06499_ _06500_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux4_1
XFILLER_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18938_ registers\[52\]\[16\] registers\[53\]\[16\] registers\[54\]\[16\] registers\[55\]\[16\]
+ _05683_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__mux4_1
.ends

