magic
tech sky130A
magscale 1 2
timestamp 1762446510
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 566 824 138906 137760
<< metal2 >>
rect 3698 139200 3754 140000
rect 9218 139200 9274 140000
rect 14738 139200 14794 140000
rect 20258 139200 20314 140000
rect 25778 139200 25834 140000
rect 31298 139200 31354 140000
rect 36818 139200 36874 140000
rect 42338 139200 42394 140000
rect 47858 139200 47914 140000
rect 53378 139200 53434 140000
rect 58898 139200 58954 140000
rect 64418 139200 64474 140000
rect 69938 139200 69994 140000
rect 75458 139200 75514 140000
rect 80978 139200 81034 140000
rect 86498 139200 86554 140000
rect 92018 139200 92074 140000
rect 97538 139200 97594 140000
rect 103058 139200 103114 140000
rect 108578 139200 108634 140000
rect 114098 139200 114154 140000
rect 119618 139200 119674 140000
rect 125138 139200 125194 140000
rect 130658 139200 130714 140000
rect 136178 139200 136234 140000
rect 5722 0 5778 800
rect 6734 0 6790 800
rect 7746 0 7802 800
rect 8758 0 8814 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11794 0 11850 800
rect 12806 0 12862 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17866 0 17922 800
rect 18878 0 18934 800
rect 19890 0 19946 800
rect 20902 0 20958 800
rect 21914 0 21970 800
rect 22926 0 22982 800
rect 23938 0 23994 800
rect 24950 0 25006 800
rect 25962 0 26018 800
rect 26974 0 27030 800
rect 27986 0 28042 800
rect 28998 0 29054 800
rect 30010 0 30066 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 33046 0 33102 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39118 0 39174 800
rect 40130 0 40186 800
rect 41142 0 41198 800
rect 42154 0 42210 800
rect 43166 0 43222 800
rect 44178 0 44234 800
rect 45190 0 45246 800
rect 46202 0 46258 800
rect 47214 0 47270 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52274 0 52330 800
rect 53286 0 53342 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56322 0 56378 800
rect 57334 0 57390 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60370 0 60426 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68466 0 68522 800
rect 69478 0 69534 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72514 0 72570 800
rect 73526 0 73582 800
rect 74538 0 74594 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77574 0 77630 800
rect 78586 0 78642 800
rect 79598 0 79654 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85670 0 85726 800
rect 86682 0 86738 800
rect 87694 0 87750 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90730 0 90786 800
rect 91742 0 91798 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94778 0 94834 800
rect 95790 0 95846 800
rect 96802 0 96858 800
rect 97814 0 97870 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103886 0 103942 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 107934 0 107990 800
rect 108946 0 109002 800
rect 109958 0 110014 800
rect 110970 0 111026 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 114006 0 114062 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 117042 0 117098 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121090 0 121146 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124126 0 124182 800
rect 125138 0 125194 800
rect 126150 0 126206 800
rect 127162 0 127218 800
rect 128174 0 128230 800
rect 129186 0 129242 800
rect 130198 0 130254 800
rect 131210 0 131266 800
rect 132222 0 132278 800
rect 133234 0 133290 800
rect 134246 0 134302 800
<< obsm2 >>
rect 110 139144 3642 139346
rect 3810 139144 9162 139346
rect 9330 139144 14682 139346
rect 14850 139144 20202 139346
rect 20370 139144 25722 139346
rect 25890 139144 31242 139346
rect 31410 139144 36762 139346
rect 36930 139144 42282 139346
rect 42450 139144 47802 139346
rect 47970 139144 53322 139346
rect 53490 139144 58842 139346
rect 59010 139144 64362 139346
rect 64530 139144 69882 139346
rect 70050 139144 75402 139346
rect 75570 139144 80922 139346
rect 81090 139144 86442 139346
rect 86610 139144 91962 139346
rect 92130 139144 97482 139346
rect 97650 139144 103002 139346
rect 103170 139144 108522 139346
rect 108690 139144 114042 139346
rect 114210 139144 119562 139346
rect 119730 139144 125082 139346
rect 125250 139144 130602 139346
rect 130770 139144 136122 139346
rect 136290 139144 138900 139346
rect 110 856 138900 139144
rect 110 734 5666 856
rect 5834 734 6678 856
rect 6846 734 7690 856
rect 7858 734 8702 856
rect 8870 734 9714 856
rect 9882 734 10726 856
rect 10894 734 11738 856
rect 11906 734 12750 856
rect 12918 734 13762 856
rect 13930 734 14774 856
rect 14942 734 15786 856
rect 15954 734 16798 856
rect 16966 734 17810 856
rect 17978 734 18822 856
rect 18990 734 19834 856
rect 20002 734 20846 856
rect 21014 734 21858 856
rect 22026 734 22870 856
rect 23038 734 23882 856
rect 24050 734 24894 856
rect 25062 734 25906 856
rect 26074 734 26918 856
rect 27086 734 27930 856
rect 28098 734 28942 856
rect 29110 734 29954 856
rect 30122 734 30966 856
rect 31134 734 31978 856
rect 32146 734 32990 856
rect 33158 734 34002 856
rect 34170 734 35014 856
rect 35182 734 36026 856
rect 36194 734 37038 856
rect 37206 734 38050 856
rect 38218 734 39062 856
rect 39230 734 40074 856
rect 40242 734 41086 856
rect 41254 734 42098 856
rect 42266 734 43110 856
rect 43278 734 44122 856
rect 44290 734 45134 856
rect 45302 734 46146 856
rect 46314 734 47158 856
rect 47326 734 48170 856
rect 48338 734 49182 856
rect 49350 734 50194 856
rect 50362 734 51206 856
rect 51374 734 52218 856
rect 52386 734 53230 856
rect 53398 734 54242 856
rect 54410 734 55254 856
rect 55422 734 56266 856
rect 56434 734 57278 856
rect 57446 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60314 856
rect 60482 734 61326 856
rect 61494 734 62338 856
rect 62506 734 63350 856
rect 63518 734 64362 856
rect 64530 734 65374 856
rect 65542 734 66386 856
rect 66554 734 67398 856
rect 67566 734 68410 856
rect 68578 734 69422 856
rect 69590 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72458 856
rect 72626 734 73470 856
rect 73638 734 74482 856
rect 74650 734 75494 856
rect 75662 734 76506 856
rect 76674 734 77518 856
rect 77686 734 78530 856
rect 78698 734 79542 856
rect 79710 734 80554 856
rect 80722 734 81566 856
rect 81734 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84602 856
rect 84770 734 85614 856
rect 85782 734 86626 856
rect 86794 734 87638 856
rect 87806 734 88650 856
rect 88818 734 89662 856
rect 89830 734 90674 856
rect 90842 734 91686 856
rect 91854 734 92698 856
rect 92866 734 93710 856
rect 93878 734 94722 856
rect 94890 734 95734 856
rect 95902 734 96746 856
rect 96914 734 97758 856
rect 97926 734 98770 856
rect 98938 734 99782 856
rect 99950 734 100794 856
rect 100962 734 101806 856
rect 101974 734 102818 856
rect 102986 734 103830 856
rect 103998 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106866 856
rect 107034 734 107878 856
rect 108046 734 108890 856
rect 109058 734 109902 856
rect 110070 734 110914 856
rect 111082 734 111926 856
rect 112094 734 112938 856
rect 113106 734 113950 856
rect 114118 734 114962 856
rect 115130 734 115974 856
rect 116142 734 116986 856
rect 117154 734 117998 856
rect 118166 734 119010 856
rect 119178 734 120022 856
rect 120190 734 121034 856
rect 121202 734 122046 856
rect 122214 734 123058 856
rect 123226 734 124070 856
rect 124238 734 125082 856
rect 125250 734 126094 856
rect 126262 734 127106 856
rect 127274 734 128118 856
rect 128286 734 129130 856
rect 129298 734 130142 856
rect 130310 734 131154 856
rect 131322 734 132166 856
rect 132334 734 133178 856
rect 133346 734 134190 856
rect 134358 734 138900 856
<< metal3 >>
rect 0 130840 800 130960
rect 0 129888 800 130008
rect 0 128936 800 129056
rect 0 127984 800 128104
rect 0 127032 800 127152
rect 0 126080 800 126200
rect 0 125128 800 125248
rect 0 124176 800 124296
rect 0 123224 800 123344
rect 0 122272 800 122392
rect 0 121320 800 121440
rect 0 120368 800 120488
rect 0 119416 800 119536
rect 0 118464 800 118584
rect 0 117512 800 117632
rect 0 116560 800 116680
rect 0 115608 800 115728
rect 0 114656 800 114776
rect 0 113704 800 113824
rect 0 112752 800 112872
rect 0 111800 800 111920
rect 0 110848 800 110968
rect 0 109896 800 110016
rect 0 108944 800 109064
rect 0 107992 800 108112
rect 0 107040 800 107160
rect 0 106088 800 106208
rect 0 105136 800 105256
rect 0 104184 800 104304
rect 0 103232 800 103352
rect 0 102280 800 102400
rect 0 101328 800 101448
rect 0 100376 800 100496
rect 0 99424 800 99544
rect 0 98472 800 98592
rect 0 97520 800 97640
rect 0 96568 800 96688
rect 0 95616 800 95736
rect 0 94664 800 94784
rect 0 93712 800 93832
rect 0 92760 800 92880
rect 0 91808 800 91928
rect 0 90856 800 90976
rect 0 89904 800 90024
rect 0 88952 800 89072
rect 0 88000 800 88120
rect 0 87048 800 87168
rect 0 86096 800 86216
rect 0 85144 800 85264
rect 0 84192 800 84312
rect 0 83240 800 83360
rect 0 82288 800 82408
rect 0 81336 800 81456
rect 0 80384 800 80504
rect 0 79432 800 79552
rect 0 78480 800 78600
rect 0 77528 800 77648
rect 0 76576 800 76696
rect 0 75624 800 75744
rect 0 74672 800 74792
rect 0 73720 800 73840
rect 0 72768 800 72888
rect 0 71816 800 71936
rect 0 70864 800 70984
rect 0 69912 800 70032
rect 0 68960 800 69080
rect 0 68008 800 68128
rect 0 67056 800 67176
rect 0 66104 800 66224
rect 0 65152 800 65272
rect 0 64200 800 64320
rect 0 63248 800 63368
rect 0 62296 800 62416
rect 0 61344 800 61464
rect 0 60392 800 60512
rect 0 59440 800 59560
rect 0 58488 800 58608
rect 0 57536 800 57656
rect 0 56584 800 56704
rect 0 55632 800 55752
rect 0 54680 800 54800
rect 0 53728 800 53848
rect 0 52776 800 52896
rect 0 51824 800 51944
rect 0 50872 800 50992
rect 0 49920 800 50040
rect 0 48968 800 49088
rect 0 48016 800 48136
rect 0 47064 800 47184
rect 0 46112 800 46232
rect 0 45160 800 45280
rect 0 44208 800 44328
rect 0 43256 800 43376
rect 0 42304 800 42424
rect 0 41352 800 41472
rect 0 40400 800 40520
rect 0 39448 800 39568
rect 0 38496 800 38616
rect 0 37544 800 37664
rect 0 36592 800 36712
rect 0 35640 800 35760
rect 0 34688 800 34808
rect 0 33736 800 33856
rect 0 32784 800 32904
rect 0 31832 800 31952
rect 0 30880 800 31000
rect 0 29928 800 30048
rect 0 28976 800 29096
rect 0 28024 800 28144
rect 0 27072 800 27192
rect 0 26120 800 26240
rect 0 25168 800 25288
rect 0 24216 800 24336
rect 0 23264 800 23384
rect 0 22312 800 22432
rect 0 21360 800 21480
rect 0 20408 800 20528
rect 0 19456 800 19576
rect 0 18504 800 18624
rect 0 17552 800 17672
rect 0 16600 800 16720
rect 0 15648 800 15768
rect 0 14696 800 14816
rect 0 13744 800 13864
rect 0 12792 800 12912
rect 0 11840 800 11960
rect 0 10888 800 11008
rect 0 9936 800 10056
rect 0 8984 800 9104
<< obsm3 >>
rect 105 131040 138539 137665
rect 880 130760 138539 131040
rect 105 130088 138539 130760
rect 880 129808 138539 130088
rect 105 129136 138539 129808
rect 880 128856 138539 129136
rect 105 128184 138539 128856
rect 880 127904 138539 128184
rect 105 127232 138539 127904
rect 880 126952 138539 127232
rect 105 126280 138539 126952
rect 880 126000 138539 126280
rect 105 125328 138539 126000
rect 880 125048 138539 125328
rect 105 124376 138539 125048
rect 880 124096 138539 124376
rect 105 123424 138539 124096
rect 880 123144 138539 123424
rect 105 122472 138539 123144
rect 880 122192 138539 122472
rect 105 121520 138539 122192
rect 880 121240 138539 121520
rect 105 120568 138539 121240
rect 880 120288 138539 120568
rect 105 119616 138539 120288
rect 880 119336 138539 119616
rect 105 118664 138539 119336
rect 880 118384 138539 118664
rect 105 117712 138539 118384
rect 880 117432 138539 117712
rect 105 116760 138539 117432
rect 880 116480 138539 116760
rect 105 115808 138539 116480
rect 880 115528 138539 115808
rect 105 114856 138539 115528
rect 880 114576 138539 114856
rect 105 113904 138539 114576
rect 880 113624 138539 113904
rect 105 112952 138539 113624
rect 880 112672 138539 112952
rect 105 112000 138539 112672
rect 880 111720 138539 112000
rect 105 111048 138539 111720
rect 880 110768 138539 111048
rect 105 110096 138539 110768
rect 880 109816 138539 110096
rect 105 109144 138539 109816
rect 880 108864 138539 109144
rect 105 108192 138539 108864
rect 880 107912 138539 108192
rect 105 107240 138539 107912
rect 880 106960 138539 107240
rect 105 106288 138539 106960
rect 880 106008 138539 106288
rect 105 105336 138539 106008
rect 880 105056 138539 105336
rect 105 104384 138539 105056
rect 880 104104 138539 104384
rect 105 103432 138539 104104
rect 880 103152 138539 103432
rect 105 102480 138539 103152
rect 880 102200 138539 102480
rect 105 101528 138539 102200
rect 880 101248 138539 101528
rect 105 100576 138539 101248
rect 880 100296 138539 100576
rect 105 99624 138539 100296
rect 880 99344 138539 99624
rect 105 98672 138539 99344
rect 880 98392 138539 98672
rect 105 97720 138539 98392
rect 880 97440 138539 97720
rect 105 96768 138539 97440
rect 880 96488 138539 96768
rect 105 95816 138539 96488
rect 880 95536 138539 95816
rect 105 94864 138539 95536
rect 880 94584 138539 94864
rect 105 93912 138539 94584
rect 880 93632 138539 93912
rect 105 92960 138539 93632
rect 880 92680 138539 92960
rect 105 92008 138539 92680
rect 880 91728 138539 92008
rect 105 91056 138539 91728
rect 880 90776 138539 91056
rect 105 90104 138539 90776
rect 880 89824 138539 90104
rect 105 89152 138539 89824
rect 880 88872 138539 89152
rect 105 88200 138539 88872
rect 880 87920 138539 88200
rect 105 87248 138539 87920
rect 880 86968 138539 87248
rect 105 86296 138539 86968
rect 880 86016 138539 86296
rect 105 85344 138539 86016
rect 880 85064 138539 85344
rect 105 84392 138539 85064
rect 880 84112 138539 84392
rect 105 83440 138539 84112
rect 880 83160 138539 83440
rect 105 82488 138539 83160
rect 880 82208 138539 82488
rect 105 81536 138539 82208
rect 880 81256 138539 81536
rect 105 80584 138539 81256
rect 880 80304 138539 80584
rect 105 79632 138539 80304
rect 880 79352 138539 79632
rect 105 78680 138539 79352
rect 880 78400 138539 78680
rect 105 77728 138539 78400
rect 880 77448 138539 77728
rect 105 76776 138539 77448
rect 880 76496 138539 76776
rect 105 75824 138539 76496
rect 880 75544 138539 75824
rect 105 74872 138539 75544
rect 880 74592 138539 74872
rect 105 73920 138539 74592
rect 880 73640 138539 73920
rect 105 72968 138539 73640
rect 880 72688 138539 72968
rect 105 72016 138539 72688
rect 880 71736 138539 72016
rect 105 71064 138539 71736
rect 880 70784 138539 71064
rect 105 70112 138539 70784
rect 880 69832 138539 70112
rect 105 69160 138539 69832
rect 880 68880 138539 69160
rect 105 68208 138539 68880
rect 880 67928 138539 68208
rect 105 67256 138539 67928
rect 880 66976 138539 67256
rect 105 66304 138539 66976
rect 880 66024 138539 66304
rect 105 65352 138539 66024
rect 880 65072 138539 65352
rect 105 64400 138539 65072
rect 880 64120 138539 64400
rect 105 63448 138539 64120
rect 880 63168 138539 63448
rect 105 62496 138539 63168
rect 880 62216 138539 62496
rect 105 61544 138539 62216
rect 880 61264 138539 61544
rect 105 60592 138539 61264
rect 880 60312 138539 60592
rect 105 59640 138539 60312
rect 880 59360 138539 59640
rect 105 58688 138539 59360
rect 880 58408 138539 58688
rect 105 57736 138539 58408
rect 880 57456 138539 57736
rect 105 56784 138539 57456
rect 880 56504 138539 56784
rect 105 55832 138539 56504
rect 880 55552 138539 55832
rect 105 54880 138539 55552
rect 880 54600 138539 54880
rect 105 53928 138539 54600
rect 880 53648 138539 53928
rect 105 52976 138539 53648
rect 880 52696 138539 52976
rect 105 52024 138539 52696
rect 880 51744 138539 52024
rect 105 51072 138539 51744
rect 880 50792 138539 51072
rect 105 50120 138539 50792
rect 880 49840 138539 50120
rect 105 49168 138539 49840
rect 880 48888 138539 49168
rect 105 48216 138539 48888
rect 880 47936 138539 48216
rect 105 47264 138539 47936
rect 880 46984 138539 47264
rect 105 46312 138539 46984
rect 880 46032 138539 46312
rect 105 45360 138539 46032
rect 880 45080 138539 45360
rect 105 44408 138539 45080
rect 880 44128 138539 44408
rect 105 43456 138539 44128
rect 880 43176 138539 43456
rect 105 42504 138539 43176
rect 880 42224 138539 42504
rect 105 41552 138539 42224
rect 880 41272 138539 41552
rect 105 40600 138539 41272
rect 880 40320 138539 40600
rect 105 39648 138539 40320
rect 880 39368 138539 39648
rect 105 38696 138539 39368
rect 880 38416 138539 38696
rect 105 37744 138539 38416
rect 880 37464 138539 37744
rect 105 36792 138539 37464
rect 880 36512 138539 36792
rect 105 35840 138539 36512
rect 880 35560 138539 35840
rect 105 34888 138539 35560
rect 880 34608 138539 34888
rect 105 33936 138539 34608
rect 880 33656 138539 33936
rect 105 32984 138539 33656
rect 880 32704 138539 32984
rect 105 32032 138539 32704
rect 880 31752 138539 32032
rect 105 31080 138539 31752
rect 880 30800 138539 31080
rect 105 30128 138539 30800
rect 880 29848 138539 30128
rect 105 29176 138539 29848
rect 880 28896 138539 29176
rect 105 28224 138539 28896
rect 880 27944 138539 28224
rect 105 27272 138539 27944
rect 880 26992 138539 27272
rect 105 26320 138539 26992
rect 880 26040 138539 26320
rect 105 25368 138539 26040
rect 880 25088 138539 25368
rect 105 24416 138539 25088
rect 880 24136 138539 24416
rect 105 23464 138539 24136
rect 880 23184 138539 23464
rect 105 22512 138539 23184
rect 880 22232 138539 22512
rect 105 21560 138539 22232
rect 880 21280 138539 21560
rect 105 20608 138539 21280
rect 880 20328 138539 20608
rect 105 19656 138539 20328
rect 880 19376 138539 19656
rect 105 18704 138539 19376
rect 880 18424 138539 18704
rect 105 17752 138539 18424
rect 880 17472 138539 17752
rect 105 16800 138539 17472
rect 880 16520 138539 16800
rect 105 15848 138539 16520
rect 880 15568 138539 15848
rect 105 14896 138539 15568
rect 880 14616 138539 14896
rect 105 13944 138539 14616
rect 880 13664 138539 13944
rect 105 12992 138539 13664
rect 880 12712 138539 12992
rect 105 12040 138539 12712
rect 880 11760 138539 12040
rect 105 11088 138539 11760
rect 880 10808 138539 11088
rect 105 10136 138539 10808
rect 880 9856 138539 10136
rect 105 9184 138539 9856
rect 880 8904 138539 9184
rect 105 1803 138539 8904
<< metal4 >>
rect 1794 2128 2414 137680
rect 19794 2128 20414 137680
rect 37794 2128 38414 137680
rect 55794 2128 56414 137680
rect 73794 2128 74414 137680
rect 91794 2128 92414 137680
rect 109794 2128 110414 137680
rect 127794 2128 128414 137680
<< obsm4 >>
rect 795 2483 1714 137461
rect 2494 2483 19714 137461
rect 20494 2483 37714 137461
rect 38494 2483 55714 137461
rect 56494 2483 73714 137461
rect 74494 2483 91714 137461
rect 92494 2483 109714 137461
rect 110494 2483 127714 137461
rect 128494 2483 136653 137461
<< labels >>
rlabel metal3 s 0 8984 800 9104 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 D1[0]
port 2 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 D1[10]
port 3 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 D1[11]
port 4 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 D1[12]
port 5 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 D1[13]
port 6 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 D1[14]
port 7 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 D1[15]
port 8 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 D1[16]
port 9 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 D1[17]
port 10 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 D1[18]
port 11 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 D1[19]
port 12 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 D1[1]
port 13 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 D1[20]
port 14 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 D1[21]
port 15 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 D1[22]
port 16 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 D1[23]
port 17 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 D1[24]
port 18 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 D1[25]
port 19 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 D1[26]
port 20 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 D1[27]
port 21 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 D1[28]
port 22 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 D1[29]
port 23 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 D1[2]
port 24 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 D1[30]
port 25 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 D1[31]
port 26 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 D1[32]
port 27 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 D1[33]
port 28 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 D1[34]
port 29 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 D1[35]
port 30 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 D1[36]
port 31 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 D1[37]
port 32 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 D1[38]
port 33 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 D1[39]
port 34 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 D1[3]
port 35 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 D1[40]
port 36 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 D1[41]
port 37 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 D1[42]
port 38 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 D1[43]
port 39 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 D1[44]
port 40 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 D1[45]
port 41 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 D1[46]
port 42 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 D1[47]
port 43 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 D1[48]
port 44 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 D1[49]
port 45 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 D1[4]
port 46 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 D1[50]
port 47 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 D1[51]
port 48 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 D1[52]
port 49 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 D1[53]
port 50 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 D1[54]
port 51 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 D1[55]
port 52 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 D1[56]
port 53 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 D1[57]
port 54 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 D1[58]
port 55 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 D1[59]
port 56 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 D1[5]
port 57 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 D1[60]
port 58 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 D1[61]
port 59 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 D1[62]
port 60 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 D1[63]
port 61 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 D1[6]
port 62 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 D1[7]
port 63 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 D1[8]
port 64 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 D1[9]
port 65 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 D2[0]
port 66 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 D2[10]
port 67 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 D2[11]
port 68 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 D2[12]
port 69 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 D2[13]
port 70 nsew signal output
rlabel metal3 s 0 84192 800 84312 6 D2[14]
port 71 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 D2[15]
port 72 nsew signal output
rlabel metal3 s 0 86096 800 86216 6 D2[16]
port 73 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 D2[17]
port 74 nsew signal output
rlabel metal3 s 0 88000 800 88120 6 D2[18]
port 75 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 D2[19]
port 76 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 D2[1]
port 77 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 D2[20]
port 78 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 D2[21]
port 79 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 D2[22]
port 80 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 D2[23]
port 81 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 D2[24]
port 82 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 D2[25]
port 83 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 D2[26]
port 84 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 D2[27]
port 85 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 D2[28]
port 86 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 D2[29]
port 87 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 D2[2]
port 88 nsew signal output
rlabel metal3 s 0 99424 800 99544 6 D2[30]
port 89 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 D2[31]
port 90 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 D2[32]
port 91 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 D2[33]
port 92 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 D2[34]
port 93 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 D2[35]
port 94 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 D2[36]
port 95 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 D2[37]
port 96 nsew signal output
rlabel metal3 s 0 107040 800 107160 6 D2[38]
port 97 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 D2[39]
port 98 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 D2[3]
port 99 nsew signal output
rlabel metal3 s 0 108944 800 109064 6 D2[40]
port 100 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 D2[41]
port 101 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 D2[42]
port 102 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 D2[43]
port 103 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 D2[44]
port 104 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 D2[45]
port 105 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 D2[46]
port 106 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 D2[47]
port 107 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 D2[48]
port 108 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 D2[49]
port 109 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 D2[4]
port 110 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 D2[50]
port 111 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 D2[51]
port 112 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 D2[52]
port 113 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 D2[53]
port 114 nsew signal output
rlabel metal3 s 0 122272 800 122392 6 D2[54]
port 115 nsew signal output
rlabel metal3 s 0 123224 800 123344 6 D2[55]
port 116 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 D2[56]
port 117 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 D2[57]
port 118 nsew signal output
rlabel metal3 s 0 126080 800 126200 6 D2[58]
port 119 nsew signal output
rlabel metal3 s 0 127032 800 127152 6 D2[59]
port 120 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 D2[5]
port 121 nsew signal output
rlabel metal3 s 0 127984 800 128104 6 D2[60]
port 122 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 D2[61]
port 123 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 D2[62]
port 124 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 D2[63]
port 125 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 D2[6]
port 126 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 D2[7]
port 127 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 D2[8]
port 128 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 D2[9]
port 129 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 D3[0]
port 130 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 D3[10]
port 131 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 D3[11]
port 132 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 D3[12]
port 133 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 D3[13]
port 134 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 D3[14]
port 135 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 D3[15]
port 136 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 D3[16]
port 137 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 D3[17]
port 138 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 D3[18]
port 139 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 D3[19]
port 140 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 D3[1]
port 141 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 D3[20]
port 142 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 D3[21]
port 143 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 D3[22]
port 144 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 D3[23]
port 145 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 D3[24]
port 146 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 D3[25]
port 147 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 D3[26]
port 148 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 D3[27]
port 149 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 D3[28]
port 150 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 D3[29]
port 151 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 D3[2]
port 152 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 D3[30]
port 153 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 D3[31]
port 154 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 D3[32]
port 155 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 D3[33]
port 156 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 D3[34]
port 157 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 D3[35]
port 158 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 D3[36]
port 159 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 D3[37]
port 160 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 D3[38]
port 161 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 D3[39]
port 162 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 D3[3]
port 163 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 D3[40]
port 164 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 D3[41]
port 165 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 D3[42]
port 166 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 D3[43]
port 167 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 D3[44]
port 168 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 D3[45]
port 169 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 D3[46]
port 170 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 D3[47]
port 171 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 D3[48]
port 172 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 D3[49]
port 173 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 D3[4]
port 174 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 D3[50]
port 175 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 D3[51]
port 176 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 D3[52]
port 177 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 D3[53]
port 178 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 D3[54]
port 179 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 D3[55]
port 180 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 D3[56]
port 181 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 D3[57]
port 182 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 D3[58]
port 183 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 D3[59]
port 184 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 D3[5]
port 185 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 D3[60]
port 186 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 D3[61]
port 187 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 D3[62]
port 188 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 D3[63]
port 189 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 D3[6]
port 190 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 D3[7]
port 191 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 D3[8]
port 192 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 D3[9]
port 193 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 DW[0]
port 194 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 DW[10]
port 195 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 DW[11]
port 196 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 DW[12]
port 197 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 DW[13]
port 198 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 DW[14]
port 199 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 DW[15]
port 200 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 DW[16]
port 201 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 DW[17]
port 202 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 DW[18]
port 203 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 DW[19]
port 204 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 DW[1]
port 205 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 DW[20]
port 206 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 DW[21]
port 207 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 DW[22]
port 208 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 DW[23]
port 209 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 DW[24]
port 210 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 DW[25]
port 211 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 DW[26]
port 212 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 DW[27]
port 213 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 DW[28]
port 214 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 DW[29]
port 215 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 DW[2]
port 216 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 DW[30]
port 217 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 DW[31]
port 218 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 DW[32]
port 219 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 DW[33]
port 220 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 DW[34]
port 221 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 DW[35]
port 222 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 DW[36]
port 223 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 DW[37]
port 224 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 DW[38]
port 225 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 DW[39]
port 226 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 DW[3]
port 227 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 DW[40]
port 228 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 DW[41]
port 229 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 DW[42]
port 230 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 DW[43]
port 231 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 DW[44]
port 232 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 DW[45]
port 233 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 DW[46]
port 234 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 DW[47]
port 235 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 DW[48]
port 236 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 DW[49]
port 237 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 DW[4]
port 238 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 DW[50]
port 239 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 DW[51]
port 240 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 DW[52]
port 241 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 DW[53]
port 242 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 DW[54]
port 243 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 DW[55]
port 244 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 DW[56]
port 245 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 DW[57]
port 246 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 DW[58]
port 247 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 DW[59]
port 248 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 DW[5]
port 249 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 DW[60]
port 250 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 DW[61]
port 251 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 DW[62]
port 252 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 DW[63]
port 253 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 DW[6]
port 254 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 DW[7]
port 255 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 DW[8]
port 256 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 DW[9]
port 257 nsew signal input
rlabel metal2 s 9218 139200 9274 140000 6 R1[0]
port 258 nsew signal input
rlabel metal2 s 14738 139200 14794 140000 6 R1[1]
port 259 nsew signal input
rlabel metal2 s 20258 139200 20314 140000 6 R1[2]
port 260 nsew signal input
rlabel metal2 s 25778 139200 25834 140000 6 R1[3]
port 261 nsew signal input
rlabel metal2 s 31298 139200 31354 140000 6 R1[4]
port 262 nsew signal input
rlabel metal2 s 36818 139200 36874 140000 6 R1[5]
port 263 nsew signal input
rlabel metal2 s 42338 139200 42394 140000 6 R2[0]
port 264 nsew signal input
rlabel metal2 s 47858 139200 47914 140000 6 R2[1]
port 265 nsew signal input
rlabel metal2 s 53378 139200 53434 140000 6 R2[2]
port 266 nsew signal input
rlabel metal2 s 58898 139200 58954 140000 6 R2[3]
port 267 nsew signal input
rlabel metal2 s 64418 139200 64474 140000 6 R2[4]
port 268 nsew signal input
rlabel metal2 s 69938 139200 69994 140000 6 R2[5]
port 269 nsew signal input
rlabel metal2 s 75458 139200 75514 140000 6 R3[0]
port 270 nsew signal input
rlabel metal2 s 80978 139200 81034 140000 6 R3[1]
port 271 nsew signal input
rlabel metal2 s 86498 139200 86554 140000 6 R3[2]
port 272 nsew signal input
rlabel metal2 s 92018 139200 92074 140000 6 R3[3]
port 273 nsew signal input
rlabel metal2 s 97538 139200 97594 140000 6 R3[4]
port 274 nsew signal input
rlabel metal2 s 103058 139200 103114 140000 6 R3[5]
port 275 nsew signal input
rlabel metal2 s 108578 139200 108634 140000 6 RW[0]
port 276 nsew signal input
rlabel metal2 s 114098 139200 114154 140000 6 RW[1]
port 277 nsew signal input
rlabel metal2 s 119618 139200 119674 140000 6 RW[2]
port 278 nsew signal input
rlabel metal2 s 125138 139200 125194 140000 6 RW[3]
port 279 nsew signal input
rlabel metal2 s 130658 139200 130714 140000 6 RW[4]
port 280 nsew signal input
rlabel metal2 s 136178 139200 136234 140000 6 RW[5]
port 281 nsew signal input
rlabel metal4 s 19794 2128 20414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 127794 2128 128414 137680 6 VGND
port 282 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 137680 6 VPWR
port 283 nsew power bidirectional
rlabel metal2 s 3698 139200 3754 140000 6 WE
port 284 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 69514186
string GDS_FILE /home/friday/check/mpw/caravel_user_project/openlane/Microwatt_FP_DFFRFile/runs/25_11_06_21_38/results/signoff/Microwatt_FP_DFFRFile.magic.gds
string GDS_START 345330
<< end >>

