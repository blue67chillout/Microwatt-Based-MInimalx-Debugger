VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Microwatt_FP_DFFRFile
  CLASS BLOCK ;
  FOREIGN Microwatt_FP_DFFRFile ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END CLK
  PIN D1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END D1[31]
  PIN D1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END D1[32]
  PIN D1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END D1[33]
  PIN D1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END D1[34]
  PIN D1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END D1[35]
  PIN D1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END D1[36]
  PIN D1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END D1[37]
  PIN D1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END D1[38]
  PIN D1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END D1[39]
  PIN D1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END D1[3]
  PIN D1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END D1[40]
  PIN D1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END D1[41]
  PIN D1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END D1[42]
  PIN D1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END D1[43]
  PIN D1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END D1[44]
  PIN D1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END D1[45]
  PIN D1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END D1[46]
  PIN D1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END D1[47]
  PIN D1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END D1[48]
  PIN D1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END D1[49]
  PIN D1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END D1[4]
  PIN D1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END D1[50]
  PIN D1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END D1[51]
  PIN D1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END D1[52]
  PIN D1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END D1[53]
  PIN D1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END D1[54]
  PIN D1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END D1[55]
  PIN D1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END D1[56]
  PIN D1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END D1[57]
  PIN D1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END D1[58]
  PIN D1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END D1[59]
  PIN D1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END D1[5]
  PIN D1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END D1[60]
  PIN D1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END D1[61]
  PIN D1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END D1[62]
  PIN D1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END D1[63]
  PIN D1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END D2[31]
  PIN D2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END D2[32]
  PIN D2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END D2[33]
  PIN D2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END D2[34]
  PIN D2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END D2[35]
  PIN D2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END D2[36]
  PIN D2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END D2[37]
  PIN D2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END D2[38]
  PIN D2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END D2[39]
  PIN D2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END D2[3]
  PIN D2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END D2[40]
  PIN D2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END D2[41]
  PIN D2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END D2[42]
  PIN D2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END D2[43]
  PIN D2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END D2[44]
  PIN D2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END D2[45]
  PIN D2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END D2[46]
  PIN D2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END D2[47]
  PIN D2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END D2[48]
  PIN D2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END D2[49]
  PIN D2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END D2[4]
  PIN D2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END D2[50]
  PIN D2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END D2[51]
  PIN D2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END D2[52]
  PIN D2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END D2[53]
  PIN D2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END D2[54]
  PIN D2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END D2[55]
  PIN D2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END D2[56]
  PIN D2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END D2[57]
  PIN D2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END D2[58]
  PIN D2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END D2[59]
  PIN D2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END D2[5]
  PIN D2[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END D2[60]
  PIN D2[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END D2[61]
  PIN D2[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END D2[62]
  PIN D2[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END D2[63]
  PIN D2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END D2[9]
  PIN D3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END D3[0]
  PIN D3[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END D3[10]
  PIN D3[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END D3[11]
  PIN D3[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END D3[12]
  PIN D3[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END D3[13]
  PIN D3[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END D3[14]
  PIN D3[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END D3[15]
  PIN D3[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END D3[16]
  PIN D3[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END D3[17]
  PIN D3[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END D3[18]
  PIN D3[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END D3[19]
  PIN D3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END D3[1]
  PIN D3[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END D3[20]
  PIN D3[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END D3[21]
  PIN D3[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END D3[22]
  PIN D3[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END D3[23]
  PIN D3[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END D3[24]
  PIN D3[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END D3[25]
  PIN D3[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END D3[26]
  PIN D3[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END D3[27]
  PIN D3[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END D3[28]
  PIN D3[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END D3[29]
  PIN D3[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END D3[2]
  PIN D3[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END D3[30]
  PIN D3[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END D3[31]
  PIN D3[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END D3[32]
  PIN D3[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END D3[33]
  PIN D3[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END D3[34]
  PIN D3[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END D3[35]
  PIN D3[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END D3[36]
  PIN D3[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END D3[37]
  PIN D3[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END D3[38]
  PIN D3[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END D3[39]
  PIN D3[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END D3[3]
  PIN D3[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END D3[40]
  PIN D3[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END D3[41]
  PIN D3[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END D3[42]
  PIN D3[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END D3[43]
  PIN D3[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END D3[44]
  PIN D3[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END D3[45]
  PIN D3[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END D3[46]
  PIN D3[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END D3[47]
  PIN D3[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END D3[48]
  PIN D3[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END D3[49]
  PIN D3[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END D3[4]
  PIN D3[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END D3[50]
  PIN D3[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END D3[51]
  PIN D3[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END D3[52]
  PIN D3[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END D3[53]
  PIN D3[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END D3[54]
  PIN D3[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END D3[55]
  PIN D3[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END D3[56]
  PIN D3[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END D3[57]
  PIN D3[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END D3[58]
  PIN D3[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END D3[59]
  PIN D3[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END D3[5]
  PIN D3[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END D3[60]
  PIN D3[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END D3[61]
  PIN D3[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END D3[62]
  PIN D3[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END D3[63]
  PIN D3[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END D3[6]
  PIN D3[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END D3[7]
  PIN D3[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END D3[8]
  PIN D3[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END D3[9]
  PIN DW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END DW[0]
  PIN DW[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END DW[10]
  PIN DW[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END DW[11]
  PIN DW[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END DW[12]
  PIN DW[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END DW[13]
  PIN DW[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END DW[14]
  PIN DW[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END DW[15]
  PIN DW[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END DW[16]
  PIN DW[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END DW[17]
  PIN DW[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END DW[18]
  PIN DW[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END DW[19]
  PIN DW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END DW[1]
  PIN DW[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END DW[20]
  PIN DW[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END DW[21]
  PIN DW[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END DW[22]
  PIN DW[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END DW[23]
  PIN DW[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END DW[24]
  PIN DW[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END DW[25]
  PIN DW[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END DW[26]
  PIN DW[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END DW[27]
  PIN DW[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END DW[28]
  PIN DW[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END DW[29]
  PIN DW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END DW[2]
  PIN DW[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END DW[30]
  PIN DW[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END DW[31]
  PIN DW[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END DW[32]
  PIN DW[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END DW[33]
  PIN DW[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END DW[34]
  PIN DW[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END DW[35]
  PIN DW[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END DW[36]
  PIN DW[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END DW[37]
  PIN DW[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END DW[38]
  PIN DW[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END DW[39]
  PIN DW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END DW[3]
  PIN DW[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END DW[40]
  PIN DW[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END DW[41]
  PIN DW[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END DW[42]
  PIN DW[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END DW[43]
  PIN DW[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END DW[44]
  PIN DW[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END DW[45]
  PIN DW[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END DW[46]
  PIN DW[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END DW[47]
  PIN DW[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END DW[48]
  PIN DW[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END DW[49]
  PIN DW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END DW[4]
  PIN DW[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END DW[50]
  PIN DW[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END DW[51]
  PIN DW[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END DW[52]
  PIN DW[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END DW[53]
  PIN DW[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END DW[54]
  PIN DW[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END DW[55]
  PIN DW[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END DW[56]
  PIN DW[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END DW[57]
  PIN DW[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END DW[58]
  PIN DW[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END DW[59]
  PIN DW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END DW[5]
  PIN DW[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END DW[60]
  PIN DW[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END DW[61]
  PIN DW[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END DW[62]
  PIN DW[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END DW[63]
  PIN DW[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END DW[6]
  PIN DW[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END DW[7]
  PIN DW[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END DW[8]
  PIN DW[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END DW[9]
  PIN R1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 696.000 46.370 700.000 ;
    END
  END R1[0]
  PIN R1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 73.690 696.000 73.970 700.000 ;
    END
  END R1[1]
  PIN R1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 101.290 696.000 101.570 700.000 ;
    END
  END R1[2]
  PIN R1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 696.000 129.170 700.000 ;
    END
  END R1[3]
  PIN R1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 156.490 696.000 156.770 700.000 ;
    END
  END R1[4]
  PIN R1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 184.090 696.000 184.370 700.000 ;
    END
  END R1[5]
  PIN R2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 211.690 696.000 211.970 700.000 ;
    END
  END R2[0]
  PIN R2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 239.290 696.000 239.570 700.000 ;
    END
  END R2[1]
  PIN R2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 266.890 696.000 267.170 700.000 ;
    END
  END R2[2]
  PIN R2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.490 696.000 294.770 700.000 ;
    END
  END R2[3]
  PIN R2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 322.090 696.000 322.370 700.000 ;
    END
  END R2[4]
  PIN R2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 349.690 696.000 349.970 700.000 ;
    END
  END R2[5]
  PIN R3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 377.290 696.000 377.570 700.000 ;
    END
  END R3[0]
  PIN R3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 404.890 696.000 405.170 700.000 ;
    END
  END R3[1]
  PIN R3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 432.490 696.000 432.770 700.000 ;
    END
  END R3[2]
  PIN R3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 460.090 696.000 460.370 700.000 ;
    END
  END R3[3]
  PIN R3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 487.690 696.000 487.970 700.000 ;
    END
  END R3[4]
  PIN R3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 515.290 696.000 515.570 700.000 ;
    END
  END R3[5]
  PIN RW[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 542.890 696.000 543.170 700.000 ;
    END
  END RW[0]
  PIN RW[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.490 696.000 570.770 700.000 ;
    END
  END RW[1]
  PIN RW[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 598.090 696.000 598.370 700.000 ;
    END
  END RW[2]
  PIN RW[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 625.690 696.000 625.970 700.000 ;
    END
  END RW[3]
  PIN RW[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 653.290 696.000 653.570 700.000 ;
    END
  END RW[4]
  PIN RW[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 680.890 696.000 681.170 700.000 ;
    END
  END RW[5]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 27.570 10.640 30.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 10.640 210.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 10.640 390.670 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 10.640 570.670 688.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 688.400 ;
    END
  END VPWR
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 18.490 696.000 18.770 700.000 ;
    END
  END WE
  OBS
      LAYER nwell ;
        RECT 5.330 10.760 694.330 688.350 ;
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 1.450 5.140 694.440 689.820 ;
      LAYER met2 ;
        RECT 0.090 695.720 18.210 696.730 ;
        RECT 19.050 695.720 45.810 696.730 ;
        RECT 46.650 695.720 73.410 696.730 ;
        RECT 74.250 695.720 101.010 696.730 ;
        RECT 101.850 695.720 128.610 696.730 ;
        RECT 129.450 695.720 156.210 696.730 ;
        RECT 157.050 695.720 183.810 696.730 ;
        RECT 184.650 695.720 211.410 696.730 ;
        RECT 212.250 695.720 239.010 696.730 ;
        RECT 239.850 695.720 266.610 696.730 ;
        RECT 267.450 695.720 294.210 696.730 ;
        RECT 295.050 695.720 321.810 696.730 ;
        RECT 322.650 695.720 349.410 696.730 ;
        RECT 350.250 695.720 377.010 696.730 ;
        RECT 377.850 695.720 404.610 696.730 ;
        RECT 405.450 695.720 432.210 696.730 ;
        RECT 433.050 695.720 459.810 696.730 ;
        RECT 460.650 695.720 487.410 696.730 ;
        RECT 488.250 695.720 515.010 696.730 ;
        RECT 515.850 695.720 542.610 696.730 ;
        RECT 543.450 695.720 570.210 696.730 ;
        RECT 571.050 695.720 597.810 696.730 ;
        RECT 598.650 695.720 625.410 696.730 ;
        RECT 626.250 695.720 653.010 696.730 ;
        RECT 653.850 695.720 680.610 696.730 ;
        RECT 681.450 695.720 693.120 696.730 ;
        RECT 0.090 4.280 693.120 695.720 ;
        RECT 0.090 3.670 28.330 4.280 ;
        RECT 29.170 3.670 33.390 4.280 ;
        RECT 34.230 3.670 38.450 4.280 ;
        RECT 39.290 3.670 43.510 4.280 ;
        RECT 44.350 3.670 48.570 4.280 ;
        RECT 49.410 3.670 53.630 4.280 ;
        RECT 54.470 3.670 58.690 4.280 ;
        RECT 59.530 3.670 63.750 4.280 ;
        RECT 64.590 3.670 68.810 4.280 ;
        RECT 69.650 3.670 73.870 4.280 ;
        RECT 74.710 3.670 78.930 4.280 ;
        RECT 79.770 3.670 83.990 4.280 ;
        RECT 84.830 3.670 89.050 4.280 ;
        RECT 89.890 3.670 94.110 4.280 ;
        RECT 94.950 3.670 99.170 4.280 ;
        RECT 100.010 3.670 104.230 4.280 ;
        RECT 105.070 3.670 109.290 4.280 ;
        RECT 110.130 3.670 114.350 4.280 ;
        RECT 115.190 3.670 119.410 4.280 ;
        RECT 120.250 3.670 124.470 4.280 ;
        RECT 125.310 3.670 129.530 4.280 ;
        RECT 130.370 3.670 134.590 4.280 ;
        RECT 135.430 3.670 139.650 4.280 ;
        RECT 140.490 3.670 144.710 4.280 ;
        RECT 145.550 3.670 149.770 4.280 ;
        RECT 150.610 3.670 154.830 4.280 ;
        RECT 155.670 3.670 159.890 4.280 ;
        RECT 160.730 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.010 4.280 ;
        RECT 170.850 3.670 175.070 4.280 ;
        RECT 175.910 3.670 180.130 4.280 ;
        RECT 180.970 3.670 185.190 4.280 ;
        RECT 186.030 3.670 190.250 4.280 ;
        RECT 191.090 3.670 195.310 4.280 ;
        RECT 196.150 3.670 200.370 4.280 ;
        RECT 201.210 3.670 205.430 4.280 ;
        RECT 206.270 3.670 210.490 4.280 ;
        RECT 211.330 3.670 215.550 4.280 ;
        RECT 216.390 3.670 220.610 4.280 ;
        RECT 221.450 3.670 225.670 4.280 ;
        RECT 226.510 3.670 230.730 4.280 ;
        RECT 231.570 3.670 235.790 4.280 ;
        RECT 236.630 3.670 240.850 4.280 ;
        RECT 241.690 3.670 245.910 4.280 ;
        RECT 246.750 3.670 250.970 4.280 ;
        RECT 251.810 3.670 256.030 4.280 ;
        RECT 256.870 3.670 261.090 4.280 ;
        RECT 261.930 3.670 266.150 4.280 ;
        RECT 266.990 3.670 271.210 4.280 ;
        RECT 272.050 3.670 276.270 4.280 ;
        RECT 277.110 3.670 281.330 4.280 ;
        RECT 282.170 3.670 286.390 4.280 ;
        RECT 287.230 3.670 291.450 4.280 ;
        RECT 292.290 3.670 296.510 4.280 ;
        RECT 297.350 3.670 301.570 4.280 ;
        RECT 302.410 3.670 306.630 4.280 ;
        RECT 307.470 3.670 311.690 4.280 ;
        RECT 312.530 3.670 316.750 4.280 ;
        RECT 317.590 3.670 321.810 4.280 ;
        RECT 322.650 3.670 326.870 4.280 ;
        RECT 327.710 3.670 331.930 4.280 ;
        RECT 332.770 3.670 336.990 4.280 ;
        RECT 337.830 3.670 342.050 4.280 ;
        RECT 342.890 3.670 347.110 4.280 ;
        RECT 347.950 3.670 352.170 4.280 ;
        RECT 353.010 3.670 357.230 4.280 ;
        RECT 358.070 3.670 362.290 4.280 ;
        RECT 363.130 3.670 367.350 4.280 ;
        RECT 368.190 3.670 372.410 4.280 ;
        RECT 373.250 3.670 377.470 4.280 ;
        RECT 378.310 3.670 382.530 4.280 ;
        RECT 383.370 3.670 387.590 4.280 ;
        RECT 388.430 3.670 392.650 4.280 ;
        RECT 393.490 3.670 397.710 4.280 ;
        RECT 398.550 3.670 402.770 4.280 ;
        RECT 403.610 3.670 407.830 4.280 ;
        RECT 408.670 3.670 412.890 4.280 ;
        RECT 413.730 3.670 417.950 4.280 ;
        RECT 418.790 3.670 423.010 4.280 ;
        RECT 423.850 3.670 428.070 4.280 ;
        RECT 428.910 3.670 433.130 4.280 ;
        RECT 433.970 3.670 438.190 4.280 ;
        RECT 439.030 3.670 443.250 4.280 ;
        RECT 444.090 3.670 448.310 4.280 ;
        RECT 449.150 3.670 453.370 4.280 ;
        RECT 454.210 3.670 458.430 4.280 ;
        RECT 459.270 3.670 463.490 4.280 ;
        RECT 464.330 3.670 468.550 4.280 ;
        RECT 469.390 3.670 473.610 4.280 ;
        RECT 474.450 3.670 478.670 4.280 ;
        RECT 479.510 3.670 483.730 4.280 ;
        RECT 484.570 3.670 488.790 4.280 ;
        RECT 489.630 3.670 493.850 4.280 ;
        RECT 494.690 3.670 498.910 4.280 ;
        RECT 499.750 3.670 503.970 4.280 ;
        RECT 504.810 3.670 509.030 4.280 ;
        RECT 509.870 3.670 514.090 4.280 ;
        RECT 514.930 3.670 519.150 4.280 ;
        RECT 519.990 3.670 524.210 4.280 ;
        RECT 525.050 3.670 529.270 4.280 ;
        RECT 530.110 3.670 534.330 4.280 ;
        RECT 535.170 3.670 539.390 4.280 ;
        RECT 540.230 3.670 544.450 4.280 ;
        RECT 545.290 3.670 549.510 4.280 ;
        RECT 550.350 3.670 554.570 4.280 ;
        RECT 555.410 3.670 559.630 4.280 ;
        RECT 560.470 3.670 564.690 4.280 ;
        RECT 565.530 3.670 569.750 4.280 ;
        RECT 570.590 3.670 574.810 4.280 ;
        RECT 575.650 3.670 579.870 4.280 ;
        RECT 580.710 3.670 584.930 4.280 ;
        RECT 585.770 3.670 589.990 4.280 ;
        RECT 590.830 3.670 595.050 4.280 ;
        RECT 595.890 3.670 600.110 4.280 ;
        RECT 600.950 3.670 605.170 4.280 ;
        RECT 606.010 3.670 610.230 4.280 ;
        RECT 611.070 3.670 615.290 4.280 ;
        RECT 616.130 3.670 620.350 4.280 ;
        RECT 621.190 3.670 625.410 4.280 ;
        RECT 626.250 3.670 630.470 4.280 ;
        RECT 631.310 3.670 635.530 4.280 ;
        RECT 636.370 3.670 640.590 4.280 ;
        RECT 641.430 3.670 645.650 4.280 ;
        RECT 646.490 3.670 650.710 4.280 ;
        RECT 651.550 3.670 655.770 4.280 ;
        RECT 656.610 3.670 660.830 4.280 ;
        RECT 661.670 3.670 665.890 4.280 ;
        RECT 666.730 3.670 670.950 4.280 ;
        RECT 671.790 3.670 693.120 4.280 ;
      LAYER met3 ;
        RECT 0.065 611.680 692.235 688.325 ;
        RECT 4.400 610.280 692.235 611.680 ;
        RECT 0.065 607.600 692.235 610.280 ;
        RECT 4.400 606.200 692.235 607.600 ;
        RECT 0.065 603.520 692.235 606.200 ;
        RECT 4.400 602.120 692.235 603.520 ;
        RECT 0.065 599.440 692.235 602.120 ;
        RECT 4.400 598.040 692.235 599.440 ;
        RECT 0.065 595.360 692.235 598.040 ;
        RECT 4.400 593.960 692.235 595.360 ;
        RECT 0.065 591.280 692.235 593.960 ;
        RECT 4.400 589.880 692.235 591.280 ;
        RECT 0.065 587.200 692.235 589.880 ;
        RECT 4.400 585.800 692.235 587.200 ;
        RECT 0.065 583.120 692.235 585.800 ;
        RECT 4.400 581.720 692.235 583.120 ;
        RECT 0.065 579.040 692.235 581.720 ;
        RECT 4.400 577.640 692.235 579.040 ;
        RECT 0.065 574.960 692.235 577.640 ;
        RECT 4.400 573.560 692.235 574.960 ;
        RECT 0.065 570.880 692.235 573.560 ;
        RECT 4.400 569.480 692.235 570.880 ;
        RECT 0.065 566.800 692.235 569.480 ;
        RECT 4.400 565.400 692.235 566.800 ;
        RECT 0.065 562.720 692.235 565.400 ;
        RECT 4.400 561.320 692.235 562.720 ;
        RECT 0.065 558.640 692.235 561.320 ;
        RECT 4.400 557.240 692.235 558.640 ;
        RECT 0.065 554.560 692.235 557.240 ;
        RECT 4.400 553.160 692.235 554.560 ;
        RECT 0.065 550.480 692.235 553.160 ;
        RECT 4.400 549.080 692.235 550.480 ;
        RECT 0.065 546.400 692.235 549.080 ;
        RECT 4.400 545.000 692.235 546.400 ;
        RECT 0.065 542.320 692.235 545.000 ;
        RECT 4.400 540.920 692.235 542.320 ;
        RECT 0.065 538.240 692.235 540.920 ;
        RECT 4.400 536.840 692.235 538.240 ;
        RECT 0.065 534.160 692.235 536.840 ;
        RECT 4.400 532.760 692.235 534.160 ;
        RECT 0.065 530.080 692.235 532.760 ;
        RECT 4.400 528.680 692.235 530.080 ;
        RECT 0.065 526.000 692.235 528.680 ;
        RECT 4.400 524.600 692.235 526.000 ;
        RECT 0.065 521.920 692.235 524.600 ;
        RECT 4.400 520.520 692.235 521.920 ;
        RECT 0.065 517.840 692.235 520.520 ;
        RECT 4.400 516.440 692.235 517.840 ;
        RECT 0.065 513.760 692.235 516.440 ;
        RECT 4.400 512.360 692.235 513.760 ;
        RECT 0.065 509.680 692.235 512.360 ;
        RECT 4.400 508.280 692.235 509.680 ;
        RECT 0.065 505.600 692.235 508.280 ;
        RECT 4.400 504.200 692.235 505.600 ;
        RECT 0.065 501.520 692.235 504.200 ;
        RECT 4.400 500.120 692.235 501.520 ;
        RECT 0.065 497.440 692.235 500.120 ;
        RECT 4.400 496.040 692.235 497.440 ;
        RECT 0.065 493.360 692.235 496.040 ;
        RECT 4.400 491.960 692.235 493.360 ;
        RECT 0.065 489.280 692.235 491.960 ;
        RECT 4.400 487.880 692.235 489.280 ;
        RECT 0.065 485.200 692.235 487.880 ;
        RECT 4.400 483.800 692.235 485.200 ;
        RECT 0.065 481.120 692.235 483.800 ;
        RECT 4.400 479.720 692.235 481.120 ;
        RECT 0.065 477.040 692.235 479.720 ;
        RECT 4.400 475.640 692.235 477.040 ;
        RECT 0.065 472.960 692.235 475.640 ;
        RECT 4.400 471.560 692.235 472.960 ;
        RECT 0.065 468.880 692.235 471.560 ;
        RECT 4.400 467.480 692.235 468.880 ;
        RECT 0.065 464.800 692.235 467.480 ;
        RECT 4.400 463.400 692.235 464.800 ;
        RECT 0.065 460.720 692.235 463.400 ;
        RECT 4.400 459.320 692.235 460.720 ;
        RECT 0.065 456.640 692.235 459.320 ;
        RECT 4.400 455.240 692.235 456.640 ;
        RECT 0.065 452.560 692.235 455.240 ;
        RECT 4.400 451.160 692.235 452.560 ;
        RECT 0.065 448.480 692.235 451.160 ;
        RECT 4.400 447.080 692.235 448.480 ;
        RECT 0.065 444.400 692.235 447.080 ;
        RECT 4.400 443.000 692.235 444.400 ;
        RECT 0.065 440.320 692.235 443.000 ;
        RECT 4.400 438.920 692.235 440.320 ;
        RECT 0.065 436.240 692.235 438.920 ;
        RECT 4.400 434.840 692.235 436.240 ;
        RECT 0.065 432.160 692.235 434.840 ;
        RECT 4.400 430.760 692.235 432.160 ;
        RECT 0.065 428.080 692.235 430.760 ;
        RECT 4.400 426.680 692.235 428.080 ;
        RECT 0.065 424.000 692.235 426.680 ;
        RECT 4.400 422.600 692.235 424.000 ;
        RECT 0.065 419.920 692.235 422.600 ;
        RECT 4.400 418.520 692.235 419.920 ;
        RECT 0.065 415.840 692.235 418.520 ;
        RECT 4.400 414.440 692.235 415.840 ;
        RECT 0.065 411.760 692.235 414.440 ;
        RECT 4.400 410.360 692.235 411.760 ;
        RECT 0.065 407.680 692.235 410.360 ;
        RECT 4.400 406.280 692.235 407.680 ;
        RECT 0.065 403.600 692.235 406.280 ;
        RECT 4.400 402.200 692.235 403.600 ;
        RECT 0.065 399.520 692.235 402.200 ;
        RECT 4.400 398.120 692.235 399.520 ;
        RECT 0.065 395.440 692.235 398.120 ;
        RECT 4.400 394.040 692.235 395.440 ;
        RECT 0.065 391.360 692.235 394.040 ;
        RECT 4.400 389.960 692.235 391.360 ;
        RECT 0.065 387.280 692.235 389.960 ;
        RECT 4.400 385.880 692.235 387.280 ;
        RECT 0.065 383.200 692.235 385.880 ;
        RECT 4.400 381.800 692.235 383.200 ;
        RECT 0.065 379.120 692.235 381.800 ;
        RECT 4.400 377.720 692.235 379.120 ;
        RECT 0.065 375.040 692.235 377.720 ;
        RECT 4.400 373.640 692.235 375.040 ;
        RECT 0.065 370.960 692.235 373.640 ;
        RECT 4.400 369.560 692.235 370.960 ;
        RECT 0.065 366.880 692.235 369.560 ;
        RECT 4.400 365.480 692.235 366.880 ;
        RECT 0.065 362.800 692.235 365.480 ;
        RECT 4.400 361.400 692.235 362.800 ;
        RECT 0.065 358.720 692.235 361.400 ;
        RECT 4.400 357.320 692.235 358.720 ;
        RECT 0.065 354.640 692.235 357.320 ;
        RECT 4.400 353.240 692.235 354.640 ;
        RECT 0.065 350.560 692.235 353.240 ;
        RECT 4.400 349.160 692.235 350.560 ;
        RECT 0.065 346.480 692.235 349.160 ;
        RECT 4.400 345.080 692.235 346.480 ;
        RECT 0.065 342.400 692.235 345.080 ;
        RECT 4.400 341.000 692.235 342.400 ;
        RECT 0.065 338.320 692.235 341.000 ;
        RECT 4.400 336.920 692.235 338.320 ;
        RECT 0.065 334.240 692.235 336.920 ;
        RECT 4.400 332.840 692.235 334.240 ;
        RECT 0.065 330.160 692.235 332.840 ;
        RECT 4.400 328.760 692.235 330.160 ;
        RECT 0.065 326.080 692.235 328.760 ;
        RECT 4.400 324.680 692.235 326.080 ;
        RECT 0.065 322.000 692.235 324.680 ;
        RECT 4.400 320.600 692.235 322.000 ;
        RECT 0.065 317.920 692.235 320.600 ;
        RECT 4.400 316.520 692.235 317.920 ;
        RECT 0.065 313.840 692.235 316.520 ;
        RECT 4.400 312.440 692.235 313.840 ;
        RECT 0.065 309.760 692.235 312.440 ;
        RECT 4.400 308.360 692.235 309.760 ;
        RECT 0.065 305.680 692.235 308.360 ;
        RECT 4.400 304.280 692.235 305.680 ;
        RECT 0.065 301.600 692.235 304.280 ;
        RECT 4.400 300.200 692.235 301.600 ;
        RECT 0.065 297.520 692.235 300.200 ;
        RECT 4.400 296.120 692.235 297.520 ;
        RECT 0.065 293.440 692.235 296.120 ;
        RECT 4.400 292.040 692.235 293.440 ;
        RECT 0.065 289.360 692.235 292.040 ;
        RECT 4.400 287.960 692.235 289.360 ;
        RECT 0.065 285.280 692.235 287.960 ;
        RECT 4.400 283.880 692.235 285.280 ;
        RECT 0.065 281.200 692.235 283.880 ;
        RECT 4.400 279.800 692.235 281.200 ;
        RECT 0.065 277.120 692.235 279.800 ;
        RECT 4.400 275.720 692.235 277.120 ;
        RECT 0.065 273.040 692.235 275.720 ;
        RECT 4.400 271.640 692.235 273.040 ;
        RECT 0.065 268.960 692.235 271.640 ;
        RECT 4.400 267.560 692.235 268.960 ;
        RECT 0.065 264.880 692.235 267.560 ;
        RECT 4.400 263.480 692.235 264.880 ;
        RECT 0.065 260.800 692.235 263.480 ;
        RECT 4.400 259.400 692.235 260.800 ;
        RECT 0.065 256.720 692.235 259.400 ;
        RECT 4.400 255.320 692.235 256.720 ;
        RECT 0.065 252.640 692.235 255.320 ;
        RECT 4.400 251.240 692.235 252.640 ;
        RECT 0.065 248.560 692.235 251.240 ;
        RECT 4.400 247.160 692.235 248.560 ;
        RECT 0.065 244.480 692.235 247.160 ;
        RECT 4.400 243.080 692.235 244.480 ;
        RECT 0.065 240.400 692.235 243.080 ;
        RECT 4.400 239.000 692.235 240.400 ;
        RECT 0.065 236.320 692.235 239.000 ;
        RECT 4.400 234.920 692.235 236.320 ;
        RECT 0.065 232.240 692.235 234.920 ;
        RECT 4.400 230.840 692.235 232.240 ;
        RECT 0.065 228.160 692.235 230.840 ;
        RECT 4.400 226.760 692.235 228.160 ;
        RECT 0.065 224.080 692.235 226.760 ;
        RECT 4.400 222.680 692.235 224.080 ;
        RECT 0.065 220.000 692.235 222.680 ;
        RECT 4.400 218.600 692.235 220.000 ;
        RECT 0.065 215.920 692.235 218.600 ;
        RECT 4.400 214.520 692.235 215.920 ;
        RECT 0.065 211.840 692.235 214.520 ;
        RECT 4.400 210.440 692.235 211.840 ;
        RECT 0.065 207.760 692.235 210.440 ;
        RECT 4.400 206.360 692.235 207.760 ;
        RECT 0.065 203.680 692.235 206.360 ;
        RECT 4.400 202.280 692.235 203.680 ;
        RECT 0.065 199.600 692.235 202.280 ;
        RECT 4.400 198.200 692.235 199.600 ;
        RECT 0.065 195.520 692.235 198.200 ;
        RECT 4.400 194.120 692.235 195.520 ;
        RECT 0.065 191.440 692.235 194.120 ;
        RECT 4.400 190.040 692.235 191.440 ;
        RECT 0.065 187.360 692.235 190.040 ;
        RECT 4.400 185.960 692.235 187.360 ;
        RECT 0.065 183.280 692.235 185.960 ;
        RECT 4.400 181.880 692.235 183.280 ;
        RECT 0.065 179.200 692.235 181.880 ;
        RECT 4.400 177.800 692.235 179.200 ;
        RECT 0.065 175.120 692.235 177.800 ;
        RECT 4.400 173.720 692.235 175.120 ;
        RECT 0.065 171.040 692.235 173.720 ;
        RECT 4.400 169.640 692.235 171.040 ;
        RECT 0.065 166.960 692.235 169.640 ;
        RECT 4.400 165.560 692.235 166.960 ;
        RECT 0.065 162.880 692.235 165.560 ;
        RECT 4.400 161.480 692.235 162.880 ;
        RECT 0.065 158.800 692.235 161.480 ;
        RECT 4.400 157.400 692.235 158.800 ;
        RECT 0.065 154.720 692.235 157.400 ;
        RECT 4.400 153.320 692.235 154.720 ;
        RECT 0.065 150.640 692.235 153.320 ;
        RECT 4.400 149.240 692.235 150.640 ;
        RECT 0.065 146.560 692.235 149.240 ;
        RECT 4.400 145.160 692.235 146.560 ;
        RECT 0.065 142.480 692.235 145.160 ;
        RECT 4.400 141.080 692.235 142.480 ;
        RECT 0.065 138.400 692.235 141.080 ;
        RECT 4.400 137.000 692.235 138.400 ;
        RECT 0.065 134.320 692.235 137.000 ;
        RECT 4.400 132.920 692.235 134.320 ;
        RECT 0.065 130.240 692.235 132.920 ;
        RECT 4.400 128.840 692.235 130.240 ;
        RECT 0.065 126.160 692.235 128.840 ;
        RECT 4.400 124.760 692.235 126.160 ;
        RECT 0.065 122.080 692.235 124.760 ;
        RECT 4.400 120.680 692.235 122.080 ;
        RECT 0.065 118.000 692.235 120.680 ;
        RECT 4.400 116.600 692.235 118.000 ;
        RECT 0.065 113.920 692.235 116.600 ;
        RECT 4.400 112.520 692.235 113.920 ;
        RECT 0.065 109.840 692.235 112.520 ;
        RECT 4.400 108.440 692.235 109.840 ;
        RECT 0.065 105.760 692.235 108.440 ;
        RECT 4.400 104.360 692.235 105.760 ;
        RECT 0.065 101.680 692.235 104.360 ;
        RECT 4.400 100.280 692.235 101.680 ;
        RECT 0.065 97.600 692.235 100.280 ;
        RECT 4.400 96.200 692.235 97.600 ;
        RECT 0.065 93.520 692.235 96.200 ;
        RECT 4.400 92.120 692.235 93.520 ;
        RECT 0.065 89.440 692.235 92.120 ;
        RECT 4.400 88.040 692.235 89.440 ;
        RECT 0.065 4.255 692.235 88.040 ;
      LAYER met4 ;
        RECT 3.055 10.240 8.570 686.625 ;
        RECT 12.470 10.240 27.170 686.625 ;
        RECT 31.070 10.240 188.570 686.625 ;
        RECT 192.470 10.240 207.170 686.625 ;
        RECT 211.070 10.240 368.570 686.625 ;
        RECT 372.470 10.240 387.170 686.625 ;
        RECT 391.070 10.240 548.570 686.625 ;
        RECT 552.470 10.240 567.170 686.625 ;
        RECT 571.070 10.240 683.265 686.625 ;
        RECT 3.055 4.935 683.265 10.240 ;
  END
END Microwatt_FP_DFFRFile
END LIBRARY

